
#******
# Preview export LEF
#
#	 Preview sub-version 5.10.41_USR1.7.43
#
# TECH LIB NAME: dje_tmp_lefImport
# TECH FILE NAME: techfile.cds
#******

VERSION 5.4 ;

NAMESCASESENSITIVE ON ;

DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

UNITS
    DATABASE MICRONS 100  ;
END UNITS

 MANUFACTURINGGRID    0.060000 ;
LAYER nwell
    TYPE MASTERSLICE ;
END nwell

LAYER nactive
    TYPE MASTERSLICE ;
END nactive

LAYER pactive
    TYPE MASTERSLICE ;
END pactive

LAYER poly
    TYPE MASTERSLICE ;
END poly

LAYER glass
    TYPE MASTERSLICE ;
END glass

LAYER pad
    TYPE MASTERSLICE ;
END pad

LAYER sblock
    TYPE MASTERSLICE ;
END sblock

LAYER text
    TYPE MASTERSLICE ;
END text

LAYER res_id
    TYPE MASTERSLICE ;
END res_id

LAYER cap_id
    TYPE MASTERSLICE ;
END cap_id

LAYER metalcap
    TYPE MASTERSLICE ;
END metalcap

LAYER nodrc
    TYPE MASTERSLICE ;
END nodrc

LAYER cc
    TYPE CUT ;
    SPACING 0.48 ;
END cc

LAYER metal1
    TYPE ROUTING ;
    WIDTH 0.36 ;
    SPACING 0.36 ;
    OFFSET 0.00 ;
    PITCH 1.08 ;
    DIRECTION HORIZONTAL ;
    RESISTANCE RPERSQ 0.06000000 ;
END metal1

LAYER via
    TYPE CUT ;
    SPACING 0.36 ;
END via

LAYER metal2
    TYPE ROUTING ;
    WIDTH 0.36 ;
    SPACING 0.48 ;
    OFFSET 0.00 ;
    PITCH 1.08 ;
    DIRECTION VERTICAL ;
    RESISTANCE RPERSQ 0.08000000 ;
END metal2

LAYER via2
    TYPE CUT ;
    SPACING 0.36 ;
END via2

LAYER metal3
    TYPE ROUTING ;
    WIDTH 0.36 ;
    SPACING 0.48 ;
    OFFSET 0.00 ;
    PITCH 1.08 ;
    DIRECTION HORIZONTAL ;
    RESISTANCE RPERSQ 0.08000000 ;
END metal3

LAYER via3
    TYPE CUT ;
    SPACING 0.36 ;
END via3

LAYER metal4
    TYPE ROUTING ;
    WIDTH 0.36 ;
    SPACING 0.48 ;
    OFFSET 0.00 ;
    PITCH 1.08 ;
    DIRECTION VERTICAL ;
    RESISTANCE RPERSQ 0.08000000 ;
END metal4

LAYER via4
    TYPE CUT ;
    SPACING 0.36 ;
END via4

LAYER metal5
    TYPE ROUTING ;
    WIDTH 0.48 ;
    SPACING 0.48 ;
    OFFSET 0.00 ;
    PITCH 2.16 ;
    DIRECTION HORIZONTAL ;
    RESISTANCE RPERSQ 0.03000000 ;
END metal5

VIA M1_P
	LAYER pactive ;
	  RECT -0.24 -0.24 0.24 0.24 ;
	LAYER cc ;
	  RECT -0.12 -0.12 0.12 0.12 ;
	LAYER metal1 ;
	  RECT -0.24 -0.24 0.24 0.24 ;
END M1_P

VIA M1_N
	LAYER nactive ;
	  RECT -0.24 -0.24 0.24 0.24 ;
	LAYER cc ;
	  RECT -0.12 -0.12 0.12 0.12 ;
	LAYER metal1 ;
	  RECT -0.24 -0.24 0.24 0.24 ;
END M1_N

VIA NTAP
	LAYER nwell ;
	  RECT -0.60 -0.60 0.60 0.60 ;
	LAYER cc ;
	  RECT -0.12 -0.12 0.12 0.12 ;
	LAYER metal1 ;
	  RECT -0.24 -0.24 0.24 0.24 ;
END NTAP

VIA M1_POLY
	LAYER poly ;
	  RECT -0.24 -0.24 0.24 0.24 ;
	LAYER cc ;
	  RECT -0.12 -0.12 0.12 0.12 ;
	LAYER metal1 ;
	  RECT -0.24 -0.24 0.24 0.24 ;
END M1_POLY

VIA M2_M1 DEFAULT
    LAYER metal1 ;
        RECT -0.30 -0.30 0.30 0.30 ;
    LAYER via ;
        RECT -0.18 -0.18 0.18 0.18 ;
    LAYER metal2 ;
        RECT -0.30 -0.30 0.30 0.30 ;
END M2_M1

VIA M5_M4 DEFAULT
    LAYER metal4 ;
        RECT -0.30 -0.30 0.30 0.30 ;
    LAYER via4 ;
        RECT -0.18 -0.18 0.18 0.18 ;
    LAYER metal5 ;
        RECT -0.42 -0.42 0.42 0.42 ;
END M5_M4

VIA M4_M3 DEFAULT
    LAYER metal3 ;
        RECT -0.30 -0.30 0.30 0.30 ;
    LAYER via3 ;
        RECT -0.18 -0.18 0.18 0.18 ;
    LAYER metal4 ;
        RECT -0.30 -0.30 0.30 0.30 ;
END M4_M3

VIA M3_M2 DEFAULT
    LAYER metal2 ;
        RECT -0.30 -0.30 0.30 0.30 ;
    LAYER via2 ;
        RECT -0.18 -0.18 0.18 0.18 ;
    LAYER metal3 ;
        RECT -0.30 -0.30 0.30 0.30 ;
END M3_M2

VIARULE viagen21 GENERATE
    LAYER metal1 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.12 ;
        METALOVERHANG 0.00 ;

    LAYER metal2 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.12 ;
        METALOVERHANG 0.00 ;

    LAYER via ;
        RECT -0.18 -0.18 0.18 0.18 ;
        SPACING 0.96 BY 0.96 ;
END viagen21

VIARULE viagen54 GENERATE
    LAYER metal5 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.12 ;
        METALOVERHANG 0.00 ;

    LAYER metal4 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.12 ;
        METALOVERHANG 0.00 ;

    LAYER via4 ;
        RECT -0.18 -0.18 0.18 0.18 ;
        SPACING 1.44 BY 1.44 ;
END viagen54

VIARULE viagen43 GENERATE
    LAYER metal3 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.12 ;
        METALOVERHANG 0.00 ;

    LAYER metal4 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.12 ;
        METALOVERHANG 0.00 ;

    LAYER via3 ;
        RECT -0.18 -0.18 0.18 0.18 ;
        SPACING 0.96 BY 0.96 ;
END viagen43

VIARULE viagen32 GENERATE
    LAYER metal3 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.12 ;
        METALOVERHANG 0.00 ;

    LAYER metal2 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.12 ;
        METALOVERHANG 0.00 ;

    LAYER via2 ;
        RECT -0.18 -0.18 0.18 0.18 ;
        SPACING 0.96 BY 0.96 ;
END viagen32

VIARULE TURN1 GENERATE
    LAYER metal1 ;
        DIRECTION VERTICAL ;

    LAYER metal1 ;
        DIRECTION HORIZONTAL ;
END TURN1

VIARULE TURN2 GENERATE
    LAYER metal2 ;
        DIRECTION VERTICAL ;

    LAYER metal2 ;
        DIRECTION HORIZONTAL ;
END TURN2

VIARULE TURN3 GENERATE
    LAYER metal3 ;
        DIRECTION VERTICAL ;

    LAYER metal3 ;
        DIRECTION HORIZONTAL ;
END TURN3

VIARULE TURN4 GENERATE
    LAYER metal4 ;
        DIRECTION VERTICAL ;

    LAYER metal4 ;
        DIRECTION HORIZONTAL ;
END TURN4

VIARULE TURN5 GENERATE
    LAYER metal5 ;
        DIRECTION VERTICAL ;

    LAYER metal5 ;
        DIRECTION HORIZONTAL ;
END TURN5

SPACING
    SAMENET cc cc 0.48 STACK  ;
    SAMENET metal1 metal1 0.36 STACK  ;
    SAMENET cc via 0.00 STACK  ;
    SAMENET metal2 metal2 0.48 STACK  ;
    SAMENET via via2 0.00 STACK  ;
    SAMENET metal3 metal3 0.48 STACK  ;
    SAMENET via2 via3 0.00 STACK  ;
    SAMENET metal4 metal4 0.48 STACK  ;
    SAMENET via3 via4 0.00 STACK  ;
    SAMENET metal5 metal5 0.48 STACK  ;
    SAMENET via via 0.36 STACK  ;
    SAMENET via2 via2 0.36 STACK  ;
    SAMENET via3 via3 0.36 STACK  ;
    SAMENET via4 via4 0.36 STACK  ;
END SPACING

SITE CoreSite
    SYMMETRY Y    ;
    CLASS CORE  ;
    SIZE 1.08 BY 15.12 ;
END CoreSite

SITE IOSite
    SYMMETRY Y    ;
    CLASS PAD  ;
    SIZE 90.00 BY 300.00 ;
END IOSite

SITE CornerSite
    SYMMETRY R90    ;
    CLASS PAD  ;
    SIZE 300.00 BY 300.00 ;
END CornerSite

MACRO ABnorC
    CLASS CORE ;
    FOREIGN ABnorC 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.48 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.72 3.18 1.20 5.64 ;
        RECT  3.36 3.18 3.84 5.64 ;
        RECT  4.68 5.16 5.16 12.18 ;
        RECT  0.72 5.16 5.64 5.64 ;
        END
    END op
    PIN ip3
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  3.00 6.24 3.48 6.72 ;
        END
    END ip3
    PIN ip2
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  1.92 7.32 2.40 7.80 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 7.32 1.32 7.80 ;
        END
    END ip1
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.40 0.00 2.88 3.66 ;
        RECT  0.00 0.00 6.48 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.72 10.50 1.20 15.12 ;
        RECT  2.64 10.50 3.12 15.12 ;
        RECT  0.00 13.80 6.48 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  3.72 9.54 4.20 12.18 ;
        RECT  1.68 9.54 2.16 12.18 ;
        RECT  1.68 9.54 4.20 10.02 ;
    END
END ABnorC

MACRO ABorC
    CLASS CORE ;
    FOREIGN ABorC 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.64 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.72 3.18 7.20 12.18 ;
        RECT  6.72 6.24 7.80 6.72 ;
        END
    END op
    PIN ip3
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  3.00 6.24 3.48 6.72 ;
        END
    END ip3
    PIN ip2
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  1.92 7.32 2.40 7.80 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 7.32 1.32 7.80 ;
        END
    END ip1
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.40 0.00 2.88 3.66 ;
        RECT  5.76 0.00 6.24 3.66 ;
        RECT  0.00 0.00 8.64 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.72 10.50 1.20 15.12 ;
        RECT  2.64 10.50 3.12 15.12 ;
        RECT  5.76 10.50 6.24 15.12 ;
        RECT  0.00 13.80 8.64 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  4.68 5.16 5.16 12.18 ;
        RECT  0.72 5.16 5.64 5.64 ;
        RECT  3.36 3.18 3.84 5.64 ;
        RECT  0.72 3.18 1.20 5.64 ;
        RECT  3.72 9.54 4.20 12.18 ;
        RECT  1.68 9.54 2.16 12.18 ;
        RECT  1.68 9.54 4.20 10.02 ;
    END
END ABorC

MACRO ab_or_c_or_d
    CLASS CORE ;
    FOREIGN ab_or_c_or_d 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.72 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.40 3.00 8.88 12.36 ;
        END
    END op
    PIN ip4
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  6.24 5.16 6.72 5.64 ;
        END
    END ip4
    PIN ip3
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  4.08 7.32 4.56 7.80 ;
        END
    END ip3
    PIN ip2
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  3.00 6.24 3.48 6.72 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 5.16 1.32 5.64 ;
        END
    END ip1
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.84 0.00 1.32 3.54 ;
        RECT  4.08 0.00 4.56 3.72 ;
        RECT  6.24 0.00 6.72 3.72 ;
        RECT  7.32 0.00 7.80 3.48 ;
        RECT  0.00 0.00 9.72 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.84 10.56 1.32 15.12 ;
        RECT  3.00 10.56 3.48 15.12 ;
        RECT  7.32 10.68 7.80 15.12 ;
        RECT  0.00 13.80 9.72 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  6.24 7.32 6.72 12.24 ;
        RECT  5.16 7.32 7.74 7.80 ;
        RECT  5.16 2.88 5.64 7.80 ;
        RECT  3.00 4.08 5.64 4.56 ;
        RECT  3.00 2.88 3.48 4.56 ;
        RECT  4.08 9.48 4.56 12.24 ;
        RECT  1.92 9.48 2.40 12.24 ;
        RECT  1.92 9.48 4.56 9.96 ;
    END
END ab_or_c_or_d

MACRO and2_1
    CLASS CORE ;
    FOREIGN and2_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.40 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.08 2.94 4.56 12.36 ;
        END
    END op
    PIN ip2
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  3.00 5.16 3.48 5.64 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 7.32 1.32 7.80 ;
        END
    END ip1
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  3.00 0.00 3.48 3.42 ;
        RECT  0.00 0.00 5.40 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.84 10.68 1.32 15.12 ;
        RECT  3.00 10.68 3.48 15.12 ;
        RECT  0.00 13.80 5.40 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  1.92 6.24 2.40 12.36 ;
        RECT  0.84 6.24 3.48 6.72 ;
        RECT  0.84 2.94 1.32 6.72 ;
    END
END and2_1

MACRO and2_2
    CLASS CORE ;
    FOREIGN and2_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.40 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.08 2.76 4.56 12.36 ;
        END
    END op
    PIN ip2
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  3.00 6.24 3.48 6.72 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 7.32 1.32 7.80 ;
        END
    END ip1
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  3.00 0.00 3.48 4.44 ;
        RECT  0.00 0.00 5.40 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.84 9.00 1.32 15.12 ;
        RECT  3.00 9.00 3.48 15.12 ;
        RECT  0.00 13.80 5.40 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  1.92 6.24 2.40 12.36 ;
        RECT  1.92 7.32 3.48 7.80 ;
        RECT  0.84 6.24 2.40 6.72 ;
        RECT  0.84 2.76 1.32 6.72 ;
    END
END and2_2

MACRO and2_4
    CLASS CORE ;
    FOREIGN and2_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.48 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.08 2.76 4.56 12.36 ;
        END
    END op
    PIN ip2
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  3.00 7.32 3.48 7.80 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 7.32 1.32 7.80 ;
        END
    END ip1
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  3.00 0.00 3.48 4.44 ;
        RECT  5.16 0.00 5.64 4.44 ;
        RECT  0.00 0.00 6.48 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.84 9.00 1.32 15.12 ;
        RECT  3.00 9.00 3.48 15.12 ;
        RECT  5.16 9.00 5.64 15.12 ;
        RECT  0.00 13.80 6.48 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  1.92 6.24 2.40 12.36 ;
        RECT  0.84 6.24 3.48 6.72 ;
        RECT  0.84 2.76 1.32 6.72 ;
    END
END and2_4

MACRO and3_1
    CLASS CORE ;
    FOREIGN and3_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.48 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.16 2.94 5.64 12.36 ;
        END
    END op
    PIN ip3
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  3.00 8.40 3.48 8.88 ;
        END
    END ip3
    PIN ip2
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  1.92 5.16 2.40 5.64 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 7.32 1.32 7.80 ;
        END
    END ip1
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  4.08 0.00 4.56 3.42 ;
        RECT  0.00 0.00 6.48 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.92 10.68 2.40 15.12 ;
        RECT  4.08 10.68 4.56 15.12 ;
        RECT  0.00 13.80 6.48 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  3.00 9.84 3.48 12.36 ;
        RECT  0.84 9.84 1.32 12.36 ;
        RECT  0.84 9.84 3.48 10.32 ;
        RECT  1.92 6.24 2.40 10.32 ;
        RECT  0.84 6.24 4.56 6.72 ;
        RECT  0.84 2.94 1.32 6.72 ;
    END
END and3_1

MACRO and3_2
    CLASS CORE ;
    FOREIGN and3_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.48 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.16 2.76 5.64 12.36 ;
        END
    END op
    PIN ip3
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  4.08 6.24 4.56 6.72 ;
        END
    END ip3
    PIN ip2
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  3.00 6.24 3.48 6.72 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 6.24 1.32 6.72 ;
        END
    END ip1
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  4.08 0.00 4.56 4.44 ;
        RECT  0.00 0.00 6.48 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.92 9.00 2.40 15.12 ;
        RECT  4.08 9.00 4.56 15.12 ;
        RECT  0.00 13.80 6.48 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  3.00 7.32 3.48 12.36 ;
        RECT  0.84 7.32 1.32 12.36 ;
        RECT  3.00 7.92 4.80 8.40 ;
        RECT  0.84 7.32 3.48 7.80 ;
        RECT  1.80 5.16 2.28 7.80 ;
        RECT  0.84 5.16 2.28 5.64 ;
        RECT  0.84 2.76 1.32 5.64 ;
    END
END and3_2

MACRO and3_4
    CLASS CORE ;
    FOREIGN and3_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.56 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.86 2.76 5.34 5.64 ;
        RECT  4.86 7.32 5.34 12.36 ;
        RECT  5.16 5.16 5.64 7.80 ;
        END
    END op
    PIN ip3
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  3.00 7.32 3.48 7.80 ;
        END
    END ip3
    PIN ip2
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  1.92 5.16 2.40 5.64 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 7.32 1.32 7.80 ;
        END
    END ip1
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  3.78 0.00 4.26 4.32 ;
        RECT  6.00 0.00 6.48 4.32 ;
        RECT  0.00 0.00 7.56 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.80 9.24 2.28 15.12 ;
        RECT  3.84 9.00 4.32 15.12 ;
        RECT  5.94 9.00 6.42 15.12 ;
        RECT  0.00 13.80 7.56 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  4.02 6.18 4.62 6.78 ;
        RECT  2.82 8.40 3.30 12.36 ;
        RECT  0.78 8.40 1.26 12.36 ;
        RECT  0.78 8.40 3.30 8.88 ;
        RECT  1.80 6.24 2.28 8.88 ;
        RECT  0.78 6.18 1.38 6.78 ;
        RECT  0.78 6.24 2.28 6.72 ;
        RECT  0.84 2.76 1.32 6.78 ;
        LAYER via ;
        RECT  4.14 6.30 4.50 6.66 ;
        RECT  0.90 6.30 1.26 6.66 ;
        LAYER metal2 ;
        RECT  4.02 6.18 4.62 6.78 ;
        RECT  0.78 6.18 1.38 6.78 ;
        RECT  0.78 6.24 4.62 6.72 ;
    END
END and3_4

MACRO and4_1
    CLASS CORE ;
    FOREIGN and4_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.56 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.40 2.88 5.88 4.56 ;
        RECT  5.70 8.40 6.18 12.36 ;
        RECT  5.40 4.08 6.72 4.56 ;
        RECT  6.24 4.08 6.72 8.88 ;
        RECT  5.70 8.40 6.72 8.88 ;
        END
    END op
    PIN ip4
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  4.08 5.16 4.56 5.64 ;
        END
    END ip4
    PIN ip3
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  3.00 8.40 3.48 8.88 ;
        END
    END ip3
    PIN ip2
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  1.92 5.16 2.40 5.64 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 8.40 1.32 8.88 ;
        END
    END ip1
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  4.38 0.00 4.86 3.54 ;
        RECT  0.00 0.00 7.56 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.78 10.56 1.26 15.12 ;
        RECT  2.82 10.56 3.30 15.12 ;
        RECT  4.74 10.56 5.22 15.12 ;
        RECT  0.00 13.80 7.56 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  3.78 9.48 4.26 12.36 ;
        RECT  1.80 6.24 2.28 12.36 ;
        RECT  1.80 9.48 4.26 9.96 ;
        RECT  0.84 6.24 5.64 6.72 ;
        RECT  0.84 2.88 1.32 6.72 ;
    END
END and4_1

MACRO and4_2
    CLASS CORE ;
    FOREIGN and4_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.56 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.40 2.76 5.88 5.64 ;
        RECT  5.70 8.40 6.18 12.36 ;
        RECT  5.40 5.16 6.72 5.64 ;
        RECT  6.24 5.16 6.72 8.88 ;
        RECT  5.70 8.40 6.72 8.88 ;
        END
    END op
    PIN ip4
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  4.08 5.16 4.56 5.64 ;
        END
    END ip4
    PIN ip3
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  3.00 7.32 3.48 7.80 ;
        END
    END ip3
    PIN ip2
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  1.92 5.16 2.40 5.64 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 7.32 1.32 7.80 ;
        END
    END ip1
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  4.38 0.00 4.86 4.26 ;
        RECT  0.00 0.00 7.56 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.78 9.00 1.26 15.12 ;
        RECT  2.82 9.48 3.30 15.12 ;
        RECT  4.74 9.00 5.22 15.12 ;
        RECT  0.00 13.80 7.56 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  5.10 6.18 5.70 6.78 ;
        RECT  3.78 8.46 4.26 12.36 ;
        RECT  1.80 6.24 2.28 12.36 ;
        RECT  1.80 8.46 4.26 8.94 ;
        RECT  0.78 6.18 1.38 6.78 ;
        RECT  0.78 6.24 2.28 6.72 ;
        RECT  0.84 2.76 1.32 6.78 ;
        LAYER via ;
        RECT  5.22 6.30 5.58 6.66 ;
        RECT  0.90 6.30 1.26 6.66 ;
        LAYER metal2 ;
        RECT  5.10 6.18 5.70 6.78 ;
        RECT  0.78 6.18 1.38 6.78 ;
        RECT  0.78 6.24 5.70 6.72 ;
    END
END and4_2

MACRO and4_4
    CLASS CORE ;
    FOREIGN and4_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.56 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.40 2.76 5.88 5.64 ;
        RECT  5.70 8.40 6.18 12.36 ;
        RECT  5.40 5.16 6.72 5.64 ;
        RECT  6.24 5.16 6.72 8.88 ;
        RECT  5.70 8.40 6.72 8.88 ;
        END
    END op
    PIN ip4
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  4.08 5.16 4.56 5.64 ;
        END
    END ip4
    PIN ip3
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  3.00 7.32 3.48 7.80 ;
        END
    END ip3
    PIN ip2
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  1.92 5.16 2.40 5.64 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 7.32 1.32 7.80 ;
        END
    END ip1
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  4.38 0.00 4.86 4.26 ;
        RECT  6.48 0.00 6.96 4.26 ;
        RECT  0.00 0.00 7.56 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.78 9.24 1.26 15.12 ;
        RECT  2.82 9.24 3.30 15.12 ;
        RECT  4.74 9.24 5.22 15.12 ;
        RECT  6.66 9.24 7.14 15.12 ;
        RECT  0.00 13.80 7.56 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  5.10 6.18 5.70 6.78 ;
        RECT  3.78 8.40 4.26 12.36 ;
        RECT  1.80 6.24 2.28 12.36 ;
        RECT  1.80 8.40 4.26 8.88 ;
        RECT  0.78 6.18 1.38 6.78 ;
        RECT  0.78 6.24 2.28 6.72 ;
        RECT  0.84 2.76 1.32 6.78 ;
        LAYER via ;
        RECT  5.22 6.30 5.58 6.66 ;
        RECT  0.90 6.30 1.26 6.66 ;
        LAYER metal2 ;
        RECT  5.10 6.18 5.70 6.78 ;
        RECT  0.78 6.18 1.38 6.78 ;
        RECT  0.78 6.24 5.70 6.72 ;
    END
END and4_4

MACRO buf_1
    CLASS CORE ;
    FOREIGN buf_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.32 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.00 4.08 3.48 9.96 ;
        RECT  3.48 2.76 3.96 4.56 ;
        RECT  3.48 9.48 3.96 12.36 ;
        END
    END op
    PIN ip
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 7.32 1.32 7.80 ;
        END
    END ip
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.30 0.00 0.78 3.24 ;
        RECT  2.46 0.00 2.94 3.24 ;
        RECT  0.00 0.00 4.32 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.36 10.68 0.84 15.12 ;
        RECT  2.52 10.68 3.00 15.12 ;
        RECT  0.00 13.80 4.32 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  1.32 8.40 1.80 12.36 ;
        RECT  1.32 8.40 2.40 8.88 ;
        RECT  1.92 6.24 2.40 8.88 ;
        RECT  1.32 6.24 2.40 6.72 ;
        RECT  1.32 2.76 1.80 6.72 ;
    END
END buf_1

MACRO buf_2
    CLASS CORE ;
    FOREIGN buf_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.32 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.00 5.16 3.48 7.80 ;
        RECT  3.48 2.76 3.96 5.64 ;
        RECT  3.48 7.32 3.96 12.36 ;
        END
    END op
    PIN ip
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 7.32 1.32 7.80 ;
        END
    END ip
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.30 0.00 0.78 4.08 ;
        RECT  2.46 0.00 2.94 4.08 ;
        RECT  0.00 0.00 4.32 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.36 9.12 0.84 15.12 ;
        RECT  2.52 9.24 3.00 15.12 ;
        RECT  0.00 13.80 4.32 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  1.32 8.40 1.80 12.36 ;
        RECT  1.32 8.40 2.40 8.88 ;
        RECT  1.92 6.24 2.40 8.88 ;
        RECT  1.32 6.24 2.40 6.72 ;
        RECT  1.32 2.76 1.80 6.72 ;
    END
END buf_2

MACRO buf_4
    CLASS CORE ;
    FOREIGN buf_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.40 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.24 2.76 3.72 5.64 ;
        RECT  3.24 8.40 3.72 12.36 ;
        RECT  3.24 5.16 4.56 5.64 ;
        RECT  4.08 5.16 4.56 8.88 ;
        RECT  3.24 8.40 4.56 8.88 ;
        END
    END op
    PIN ip
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 7.32 1.32 7.80 ;
        END
    END ip
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.30 0.00 0.78 4.44 ;
        RECT  2.28 0.00 2.76 4.44 ;
        RECT  4.20 0.00 4.68 4.44 ;
        RECT  0.00 0.00 5.40 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.30 9.12 0.78 15.12 ;
        RECT  2.28 9.24 2.76 15.12 ;
        RECT  4.20 9.24 4.68 15.12 ;
        RECT  0.00 13.80 5.40 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  1.32 8.40 1.80 12.36 ;
        RECT  1.32 8.40 2.40 8.88 ;
        RECT  1.92 6.24 2.40 8.88 ;
        RECT  1.92 7.32 3.48 7.80 ;
        RECT  1.32 6.24 2.40 6.72 ;
        RECT  1.32 2.76 1.80 6.72 ;
    END
END buf_4

MACRO bufzp_2
    CLASS CORE ;
    FOREIGN bufzp_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.64 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.32 3.00 7.80 12.12 ;
        END
    END op
    PIN ip
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 7.32 1.32 7.80 ;
        END
    END ip
    PIN c
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal2 ;
        RECT  2.94 7.26 3.54 7.86 ;
        RECT  2.94 7.32 6.78 7.80 ;
        RECT  6.18 7.26 6.78 7.86 ;
        LAYER metal1 ;
        RECT  2.94 7.26 3.54 7.86 ;
        RECT  6.18 7.26 6.78 7.86 ;
        LAYER via ;
        RECT  3.06 7.38 3.42 7.74 ;
        RECT  6.30 7.38 6.66 7.74 ;
        END
    END c
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.90 0.00 1.38 3.48 ;
        RECT  3.06 0.00 3.54 3.48 ;
        RECT  5.22 0.00 5.70 4.32 ;
        RECT  0.00 0.00 8.64 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.90 10.68 1.38 15.12 ;
        RECT  3.06 10.68 3.54 15.12 ;
        RECT  5.22 9.24 5.70 15.12 ;
        RECT  0.00 13.80 8.64 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  6.18 6.18 6.78 6.78 ;
        RECT  5.10 5.10 5.70 5.70 ;
        RECT  4.08 3.00 4.56 12.36 ;
        RECT  4.02 6.18 4.62 6.78 ;
        RECT  1.92 3.00 2.40 12.36 ;
        RECT  1.86 5.10 2.46 5.70 ;
        LAYER via ;
        RECT  6.30 6.30 6.66 6.66 ;
        RECT  5.22 5.22 5.58 5.58 ;
        RECT  4.14 6.30 4.50 6.66 ;
        RECT  1.98 5.22 2.34 5.58 ;
        LAYER metal2 ;
        RECT  6.18 6.18 6.78 6.78 ;
        RECT  4.02 6.18 4.62 6.78 ;
        RECT  4.02 6.24 6.78 6.72 ;
        RECT  5.10 5.10 5.70 5.70 ;
        RECT  1.86 5.10 2.46 5.70 ;
        RECT  1.86 5.16 5.70 5.64 ;
    END
END bufzp_2

MACRO cd_12
    CLASS CORE ;
    FOREIGN cd_12 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.96 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.16 2.76 11.64 5.64 ;
        RECT  11.16 8.40 11.64 12.36 ;
        RECT  11.16 5.16 12.48 5.64 ;
        RECT  12.00 5.16 12.48 8.88 ;
        RECT  11.16 8.40 12.48 8.88 ;
        END
    END op
    PIN ip
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 7.32 1.32 7.80 ;
        END
    END ip
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.30 0.00 0.78 4.44 ;
        RECT  2.28 0.00 2.76 4.44 ;
        RECT  4.26 0.00 4.74 4.44 ;
        RECT  6.24 0.00 6.72 4.44 ;
        RECT  8.22 0.00 8.70 4.44 ;
        RECT  10.20 0.00 10.68 4.44 ;
        RECT  12.12 0.00 12.60 4.44 ;
        RECT  0.00 0.00 12.96 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.30 9.12 0.78 15.12 ;
        RECT  2.28 9.24 2.76 15.12 ;
        RECT  4.26 9.24 4.74 15.12 ;
        RECT  6.24 9.24 6.72 15.12 ;
        RECT  8.22 9.24 8.70 15.12 ;
        RECT  10.20 9.24 10.68 15.12 ;
        RECT  12.12 9.24 12.60 15.12 ;
        RECT  0.00 13.80 12.96 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  9.24 8.40 9.72 12.36 ;
        RECT  9.24 8.40 10.80 8.88 ;
        RECT  10.32 6.24 10.80 8.88 ;
        RECT  10.32 7.32 11.04 7.80 ;
        RECT  9.24 6.24 10.80 6.72 ;
        RECT  9.24 2.76 9.72 6.72 ;
        RECT  7.26 8.40 7.74 12.36 ;
        RECT  7.26 8.40 8.70 8.88 ;
        RECT  8.22 5.16 8.70 8.88 ;
        RECT  8.22 7.32 9.96 7.80 ;
        RECT  7.26 5.16 8.70 5.64 ;
        RECT  7.26 2.76 7.74 5.64 ;
        RECT  5.28 8.40 5.76 12.36 ;
        RECT  5.28 8.40 6.72 8.88 ;
        RECT  6.24 6.24 6.72 8.88 ;
        RECT  6.24 7.32 7.80 7.80 ;
        RECT  5.28 6.24 6.72 6.72 ;
        RECT  5.28 2.76 5.76 6.72 ;
        RECT  3.30 8.40 3.78 12.36 ;
        RECT  3.30 8.40 4.56 8.88 ;
        RECT  4.08 6.24 4.56 8.88 ;
        RECT  4.08 7.32 5.70 7.80 ;
        RECT  3.30 6.24 4.56 6.72 ;
        RECT  3.30 2.76 3.78 6.72 ;
        RECT  1.32 8.40 1.80 12.36 ;
        RECT  1.32 8.40 2.40 8.88 ;
        RECT  1.92 5.16 2.40 8.88 ;
        RECT  1.92 7.32 3.48 7.80 ;
        RECT  1.32 5.16 2.40 5.64 ;
        RECT  1.32 2.76 1.80 5.64 ;
    END
END cd_12

MACRO cd_16
    CLASS CORE ;
    FOREIGN cd_16 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 18.36 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  16.26 2.76 16.74 5.64 ;
        RECT  16.26 8.40 16.74 12.36 ;
        RECT  16.26 5.16 17.52 5.64 ;
        RECT  17.04 5.16 17.52 8.88 ;
        RECT  16.26 8.40 17.52 8.88 ;
        END
    END op
    PIN ip
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 7.32 1.32 7.80 ;
        END
    END ip
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.30 0.00 0.78 4.44 ;
        RECT  2.28 0.00 2.76 4.44 ;
        RECT  4.26 0.00 4.74 4.44 ;
        RECT  6.24 0.00 6.72 4.44 ;
        RECT  8.22 0.00 8.70 4.44 ;
        RECT  9.30 0.00 9.78 4.44 ;
        RECT  11.28 0.00 11.76 4.44 ;
        RECT  13.26 0.00 13.74 4.44 ;
        RECT  15.24 0.00 15.72 4.44 ;
        RECT  17.22 0.00 17.70 4.44 ;
        RECT  0.00 0.00 18.36 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.30 9.12 0.78 15.12 ;
        RECT  2.28 9.24 2.76 15.12 ;
        RECT  4.26 9.24 4.74 15.12 ;
        RECT  6.24 9.24 6.72 15.12 ;
        RECT  8.22 9.24 8.70 15.12 ;
        RECT  9.30 9.12 9.78 15.12 ;
        RECT  11.28 9.24 11.76 15.12 ;
        RECT  13.26 9.24 13.74 15.12 ;
        RECT  15.24 9.24 15.72 15.12 ;
        RECT  17.22 9.24 17.70 15.12 ;
        RECT  0.00 13.80 18.36 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  14.28 8.40 14.76 12.36 ;
        RECT  14.28 8.40 15.36 8.88 ;
        RECT  14.88 6.24 15.36 8.88 ;
        RECT  14.88 7.32 16.44 7.80 ;
        RECT  14.28 6.24 15.36 6.72 ;
        RECT  14.28 2.76 14.76 6.72 ;
        RECT  12.30 8.40 12.78 12.36 ;
        RECT  12.72 6.24 13.20 8.88 ;
        RECT  12.72 7.32 14.28 7.80 ;
        RECT  12.30 2.76 12.78 6.72 ;
        RECT  10.32 8.40 10.80 12.36 ;
        RECT  10.56 6.24 11.04 8.88 ;
        RECT  10.56 7.32 12.12 7.80 ;
        RECT  10.32 2.76 10.80 6.72 ;
        RECT  7.26 8.40 7.74 12.36 ;
        RECT  7.26 8.40 8.82 8.88 ;
        RECT  8.34 5.16 8.82 8.88 ;
        RECT  8.34 7.32 9.96 7.80 ;
        RECT  7.26 5.16 8.82 5.64 ;
        RECT  7.26 2.76 7.74 5.64 ;
        RECT  5.28 8.40 5.76 12.36 ;
        RECT  5.28 8.40 6.72 8.88 ;
        RECT  6.24 6.24 6.72 8.88 ;
        RECT  6.24 7.32 7.80 7.80 ;
        RECT  5.28 6.24 6.72 6.72 ;
        RECT  5.28 2.76 5.76 6.72 ;
        RECT  3.30 8.40 3.78 12.36 ;
        RECT  3.30 8.40 4.56 8.88 ;
        RECT  4.08 6.24 4.56 8.88 ;
        RECT  4.08 7.32 5.70 7.80 ;
        RECT  3.30 6.24 4.56 6.72 ;
        RECT  3.30 2.76 3.78 6.72 ;
        RECT  1.32 8.40 1.80 12.36 ;
        RECT  1.32 8.40 2.40 8.88 ;
        RECT  1.92 5.16 2.40 8.88 ;
        RECT  1.92 7.32 3.48 7.80 ;
        RECT  1.32 5.16 2.40 5.64 ;
        RECT  1.32 2.76 1.80 5.64 ;
    END
END cd_16

MACRO cd_8
    CLASS CORE ;
    FOREIGN cd_8 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.72 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.26 2.76 7.74 5.64 ;
        RECT  7.26 8.40 7.74 12.36 ;
        RECT  7.26 5.16 8.82 5.64 ;
        RECT  8.34 5.16 8.82 8.88 ;
        RECT  7.26 8.40 8.82 8.88 ;
        END
    END op
    PIN ip
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 7.32 1.32 7.80 ;
        END
    END ip
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.30 0.00 0.78 4.44 ;
        RECT  2.28 0.00 2.76 4.44 ;
        RECT  4.26 0.00 4.74 4.44 ;
        RECT  6.24 0.00 6.72 4.44 ;
        RECT  8.22 0.00 8.70 4.44 ;
        RECT  0.00 0.00 9.72 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.30 9.12 0.78 15.12 ;
        RECT  2.28 9.24 2.76 15.12 ;
        RECT  4.26 9.24 4.74 15.12 ;
        RECT  6.24 9.24 6.72 15.12 ;
        RECT  8.22 9.24 8.70 15.12 ;
        RECT  0.00 13.80 9.72 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  5.28 8.40 5.76 12.36 ;
        RECT  5.28 8.40 6.72 8.88 ;
        RECT  6.24 6.24 6.72 8.88 ;
        RECT  6.24 7.32 7.80 7.80 ;
        RECT  5.28 6.24 6.72 6.72 ;
        RECT  5.28 2.76 5.76 6.72 ;
        RECT  3.30 8.40 3.78 12.36 ;
        RECT  3.30 8.40 4.56 8.88 ;
        RECT  4.08 6.24 4.56 8.88 ;
        RECT  4.08 7.32 5.70 7.80 ;
        RECT  3.30 6.24 4.56 6.72 ;
        RECT  3.30 2.76 3.78 6.72 ;
        RECT  1.32 8.40 1.80 12.36 ;
        RECT  1.32 8.40 2.40 8.88 ;
        RECT  1.92 5.16 2.40 8.88 ;
        RECT  1.92 7.32 3.48 7.80 ;
        RECT  1.32 5.16 2.40 5.64 ;
        RECT  1.32 2.76 1.80 5.64 ;
    END
END cd_8

MACRO dksp_1
    CLASS CORE ;
    FOREIGN dksp_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 30.24 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN sb
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  3.00 5.10 4.20 5.70 ;
        END
    END sb
    PIN qb
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  26.70 5.10 27.72 5.70 ;
        RECT  27.24 2.76 27.72 12.36 ;
        END
    END qb
    PIN q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  28.86 6.18 29.70 6.78 ;
        RECT  29.22 2.76 29.70 12.36 ;
        END
    END q
    PIN ip
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 7.32 1.32 7.80 ;
        END
    END ip
    PIN ck
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER metal1 ;
        RECT  12.66 6.18 13.26 6.78 ;
        END
    END ck
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.66 0.00 1.14 3.60 ;
        RECT  2.64 0.00 3.12 3.60 ;
        RECT  9.18 0.00 9.66 3.60 ;
        RECT  11.16 0.00 11.64 3.60 ;
        RECT  13.14 0.00 13.62 3.60 ;
        RECT  15.12 0.00 15.60 3.60 ;
        RECT  22.26 0.00 22.74 3.60 ;
        RECT  24.24 0.00 24.72 3.60 ;
        RECT  26.22 0.00 26.70 4.44 ;
        RECT  28.20 0.00 28.68 4.44 ;
        RECT  0.00 0.00 30.24 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.66 10.68 1.14 15.12 ;
        RECT  2.64 10.68 3.12 15.12 ;
        RECT  4.68 10.68 5.16 15.12 ;
        RECT  9.18 10.68 9.66 15.12 ;
        RECT  11.16 10.68 11.64 15.12 ;
        RECT  13.14 10.68 13.62 15.12 ;
        RECT  15.12 10.68 15.60 15.12 ;
        RECT  22.26 10.68 22.74 15.12 ;
        RECT  24.24 10.68 24.72 15.12 ;
        RECT  26.22 9.00 26.70 15.12 ;
        RECT  28.20 9.00 28.68 15.12 ;
        RECT  0.00 13.80 30.24 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  28.08 7.26 28.68 7.86 ;
        RECT  25.26 2.76 25.74 12.36 ;
        RECT  25.20 7.26 25.80 7.86 ;
        RECT  23.28 2.76 23.76 12.36 ;
        RECT  23.28 4.56 24.36 5.04 ;
        RECT  22.14 6.18 22.74 6.78 ;
        RECT  20.46 7.26 20.94 12.36 ;
        RECT  20.40 7.26 21.00 7.86 ;
        RECT  20.40 7.26 21.78 7.80 ;
        RECT  21.30 3.60 21.78 7.80 ;
        RECT  20.46 3.60 21.78 4.08 ;
        RECT  20.46 2.76 20.94 4.08 ;
        RECT  20.28 4.50 20.88 5.10 ;
        RECT  19.44 2.76 19.92 12.36 ;
        RECT  20.28 6.18 20.88 6.78 ;
        RECT  19.44 6.24 20.88 6.72 ;
        RECT  18.36 5.10 18.96 5.70 ;
        RECT  18.42 7.32 18.90 12.36 ;
        RECT  18.36 8.34 18.96 8.94 ;
        RECT  17.40 7.32 18.90 7.80 ;
        RECT  17.40 3.60 17.88 7.80 ;
        RECT  17.40 3.60 18.90 4.08 ;
        RECT  18.42 2.76 18.90 4.08 ;
        RECT  17.28 9.42 17.88 10.02 ;
        RECT  16.14 2.76 16.62 12.36 ;
        RECT  16.08 5.10 16.68 5.70 ;
        RECT  14.16 2.76 14.64 12.36 ;
        RECT  14.10 9.42 14.70 10.02 ;
        RECT  14.10 7.26 14.70 7.86 ;
        RECT  14.16 6.24 15.12 6.72 ;
        RECT  14.10 4.02 14.70 4.62 ;
        RECT  12.18 7.68 12.66 12.36 ;
        RECT  12.12 9.42 12.72 10.02 ;
        RECT  11.64 7.68 12.66 8.16 ;
        RECT  11.64 4.56 12.12 8.16 ;
        RECT  11.64 4.56 12.66 5.04 ;
        RECT  12.18 2.76 12.66 5.04 ;
        RECT  10.20 2.76 10.68 12.36 ;
        RECT  10.14 8.34 10.74 8.94 ;
        RECT  10.20 6.48 11.04 6.96 ;
        RECT  9.06 8.34 9.66 8.94 ;
        RECT  8.64 5.10 9.24 5.70 ;
        RECT  8.64 7.26 9.24 7.86 ;
        RECT  7.68 2.76 8.16 12.36 ;
        RECT  7.62 9.42 8.22 10.02 ;
        RECT  6.66 2.76 7.14 12.36 ;
        RECT  6.66 8.34 7.26 8.94 ;
        RECT  5.58 4.80 6.18 5.40 ;
        RECT  5.64 7.08 6.12 12.36 ;
        RECT  3.66 7.08 4.14 12.36 ;
        RECT  3.66 7.08 6.12 7.56 ;
        RECT  4.68 2.76 5.16 7.56 ;
        RECT  5.64 2.76 6.12 4.08 ;
        RECT  4.68 2.76 6.12 3.24 ;
        RECT  1.68 2.76 2.16 12.36 ;
        LAYER via ;
        RECT  28.20 7.38 28.56 7.74 ;
        RECT  25.32 7.38 25.68 7.74 ;
        RECT  22.26 6.30 22.62 6.66 ;
        RECT  20.52 7.38 20.88 7.74 ;
        RECT  20.40 4.62 20.76 4.98 ;
        RECT  20.40 6.30 20.76 6.66 ;
        RECT  18.48 5.22 18.84 5.58 ;
        RECT  18.48 8.46 18.84 8.82 ;
        RECT  17.40 9.54 17.76 9.90 ;
        RECT  16.20 5.22 16.56 5.58 ;
        RECT  14.22 4.14 14.58 4.50 ;
        RECT  14.22 7.38 14.58 7.74 ;
        RECT  14.22 9.54 14.58 9.90 ;
        RECT  12.24 9.54 12.60 9.90 ;
        RECT  10.26 8.46 10.62 8.82 ;
        RECT  9.18 8.46 9.54 8.82 ;
        RECT  8.76 5.22 9.12 5.58 ;
        RECT  8.76 7.38 9.12 7.74 ;
        RECT  7.74 9.54 8.10 9.90 ;
        RECT  6.78 8.46 7.14 8.82 ;
        RECT  5.70 4.92 6.06 5.28 ;
        LAYER metal2 ;
        RECT  28.08 7.26 28.68 7.86 ;
        RECT  25.20 7.26 25.80 7.86 ;
        RECT  20.40 7.26 21.00 7.86 ;
        RECT  20.40 7.32 28.68 7.80 ;
        RECT  22.14 6.18 22.74 6.78 ;
        RECT  20.28 6.18 20.88 6.78 ;
        RECT  20.28 6.24 22.74 6.72 ;
        RECT  5.58 4.80 6.18 5.40 ;
        RECT  5.64 4.08 6.18 5.40 ;
        RECT  20.28 4.08 20.88 5.10 ;
        RECT  14.10 4.02 14.70 4.62 ;
        RECT  5.64 4.08 20.88 4.56 ;
        RECT  18.36 5.10 18.96 5.70 ;
        RECT  16.08 5.10 16.68 5.70 ;
        RECT  8.64 5.10 9.24 5.70 ;
        RECT  8.64 5.16 18.96 5.64 ;
        RECT  18.36 8.34 18.96 8.94 ;
        RECT  10.14 8.34 10.74 8.94 ;
        RECT  10.14 8.40 18.96 8.88 ;
        RECT  17.28 9.42 17.88 10.02 ;
        RECT  14.10 9.42 14.70 10.02 ;
        RECT  14.10 9.48 17.88 9.96 ;
        RECT  14.10 7.26 14.70 7.86 ;
        RECT  8.64 7.26 9.24 7.86 ;
        RECT  8.64 7.32 14.70 7.80 ;
        RECT  12.12 9.42 12.72 10.02 ;
        RECT  7.62 9.42 8.22 10.02 ;
        RECT  7.62 9.48 12.72 9.96 ;
        RECT  9.06 8.34 9.66 8.94 ;
        RECT  6.66 8.34 7.26 8.94 ;
        RECT  6.66 8.40 9.66 8.88 ;
    END
END dksp_1

MACRO dp_1
    CLASS CORE ;
    FOREIGN dp_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 19.44 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  17.28 8.40 17.76 12.30 ;
        RECT  15.96 6.24 18.60 6.72 ;
        RECT  18.12 4.08 18.60 8.88 ;
        RECT  17.28 8.40 18.60 8.88 ;
        RECT  18.48 2.88 18.96 4.56 ;
        END
    END q
    PIN ip
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 7.32 1.32 7.80 ;
        END
    END ip
    PIN ck
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER metal1 ;
        RECT  3.00 6.24 3.48 6.72 ;
        END
    END ck
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.30 0.00 0.78 3.48 ;
        RECT  2.46 0.00 2.94 3.48 ;
        RECT  7.86 0.00 8.34 3.48 ;
        RECT  10.38 0.00 10.86 3.48 ;
        RECT  12.48 0.00 12.96 3.48 ;
        RECT  17.34 0.00 17.82 3.48 ;
        RECT  0.00 0.00 19.44 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.30 10.62 0.78 15.12 ;
        RECT  2.46 10.62 2.94 15.12 ;
        RECT  7.50 10.62 7.98 15.12 ;
        RECT  10.38 10.62 10.86 15.12 ;
        RECT  12.48 10.62 12.96 15.12 ;
        RECT  16.26 10.62 16.74 15.12 ;
        RECT  0.00 13.80 19.44 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  14.28 9.48 14.76 12.30 ;
        RECT  13.80 7.32 14.28 9.96 ;
        RECT  13.80 7.32 17.52 7.80 ;
        RECT  14.88 4.08 15.36 7.80 ;
        RECT  14.88 4.08 15.90 4.56 ;
        RECT  15.42 2.88 15.90 4.56 ;
        RECT  15.90 5.10 16.50 5.70 ;
        RECT  14.82 8.34 15.42 8.94 ;
        RECT  13.38 3.00 14.94 3.48 ;
        RECT  13.74 6.18 14.34 6.78 ;
        RECT  13.80 4.02 14.28 6.78 ;
        RECT  13.74 4.02 14.34 4.62 ;
        RECT  11.40 9.48 11.88 12.30 ;
        RECT  11.64 4.08 12.12 9.96 ;
        RECT  11.58 7.26 12.18 7.86 ;
        RECT  11.58 7.32 13.20 7.80 ;
        RECT  11.40 2.88 11.88 4.56 ;
        RECT  5.76 7.32 6.24 12.30 ;
        RECT  5.76 8.40 10.14 8.88 ;
        RECT  9.66 7.32 10.14 8.88 ;
        RECT  9.66 7.32 11.04 7.80 ;
        RECT  5.64 2.88 6.12 7.80 ;
        RECT  8.76 2.94 9.36 3.54 ;
        RECT  7.26 4.02 7.86 4.62 ;
        RECT  7.26 7.26 7.86 7.86 ;
        RECT  6.60 2.94 7.20 3.54 ;
        RECT  4.74 10.62 5.22 12.30 ;
        RECT  4.68 11.58 5.28 12.18 ;
        RECT  4.56 2.94 5.16 3.54 ;
        RECT  3.54 9.48 4.02 12.30 ;
        RECT  3.54 9.48 4.56 9.96 ;
        RECT  4.08 4.08 4.56 9.96 ;
        RECT  4.02 6.18 4.62 6.78 ;
        RECT  3.48 4.08 4.56 4.56 ;
        RECT  3.48 2.88 3.96 4.56 ;
        RECT  2.94 8.34 3.54 8.94 ;
        RECT  1.86 4.02 2.46 4.62 ;
        RECT  1.26 2.94 1.86 3.54 ;
        RECT  1.32 10.62 1.80 12.30 ;
        RECT  1.26 11.58 1.86 12.18 ;
        LAYER via ;
        RECT  16.02 5.22 16.38 5.58 ;
        RECT  14.94 8.46 15.30 8.82 ;
        RECT  13.86 4.14 14.22 4.50 ;
        RECT  13.86 6.30 14.22 6.66 ;
        RECT  11.70 7.38 12.06 7.74 ;
        RECT  8.88 3.06 9.24 3.42 ;
        RECT  7.38 4.14 7.74 4.50 ;
        RECT  7.38 7.38 7.74 7.74 ;
        RECT  6.72 3.06 7.08 3.42 ;
        RECT  4.80 11.70 5.16 12.06 ;
        RECT  4.68 3.06 5.04 3.42 ;
        RECT  4.14 6.30 4.50 6.66 ;
        RECT  3.06 8.46 3.42 8.82 ;
        RECT  1.98 4.14 2.34 4.50 ;
        RECT  1.38 3.06 1.74 3.42 ;
        RECT  1.38 11.70 1.74 12.06 ;
        LAYER metal2 ;
        RECT  15.90 5.10 16.50 5.70 ;
        RECT  15.96 4.08 16.44 5.70 ;
        RECT  13.74 4.02 14.34 4.62 ;
        RECT  13.74 4.08 16.44 4.56 ;
        RECT  14.82 8.34 15.42 8.94 ;
        RECT  2.94 8.34 3.54 8.94 ;
        RECT  2.94 8.40 15.42 8.88 ;
        RECT  13.74 6.18 14.34 6.78 ;
        RECT  4.02 6.18 4.62 6.78 ;
        RECT  4.02 6.24 14.34 6.72 ;
        RECT  11.58 7.26 12.18 7.86 ;
        RECT  7.26 7.26 7.86 7.86 ;
        RECT  7.26 7.32 12.18 7.80 ;
        RECT  8.76 2.94 9.36 3.54 ;
        RECT  6.60 2.94 7.20 3.54 ;
        RECT  6.60 3.00 9.36 3.48 ;
        RECT  7.26 4.02 7.86 4.62 ;
        RECT  1.86 4.02 2.46 4.62 ;
        RECT  1.86 4.08 7.86 4.56 ;
        RECT  4.68 11.58 5.28 12.18 ;
        RECT  1.26 11.58 1.86 12.18 ;
        RECT  1.26 11.64 5.28 12.12 ;
        RECT  4.56 2.94 5.16 3.54 ;
        RECT  1.26 2.94 1.86 3.54 ;
        RECT  1.26 3.00 5.16 3.48 ;
    END
END dp_1

MACRO dp_2
    CLASS CORE ;
    FOREIGN dp_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 20.52 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  15.96 6.24 19.68 6.72 ;
        RECT  19.20 5.16 19.68 8.94 ;
        RECT  19.56 2.76 20.04 5.64 ;
        RECT  19.56 8.46 20.04 12.36 ;
        END
    END q
    PIN ip
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 7.32 1.32 7.80 ;
        END
    END ip
    PIN ck
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER metal1 ;
        RECT  3.00 6.24 3.48 6.72 ;
        END
    END ck
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.36 0.00 0.84 3.48 ;
        RECT  2.52 0.00 3.00 3.48 ;
        RECT  7.92 0.00 8.40 3.48 ;
        RECT  10.44 0.00 10.92 3.48 ;
        RECT  12.54 0.00 13.02 3.48 ;
        RECT  17.40 0.00 17.88 3.48 ;
        RECT  18.48 0.00 18.96 4.44 ;
        RECT  0.00 0.00 20.52 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.36 10.68 0.84 15.12 ;
        RECT  2.52 10.68 3.00 15.12 ;
        RECT  7.56 10.68 8.04 15.12 ;
        RECT  10.44 10.68 10.92 15.12 ;
        RECT  12.54 10.68 13.02 15.12 ;
        RECT  16.32 10.68 16.80 15.12 ;
        RECT  18.54 9.36 19.02 15.12 ;
        RECT  0.00 13.80 20.52 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  14.34 9.54 14.82 12.36 ;
        RECT  13.86 7.38 14.34 10.02 ;
        RECT  13.86 7.38 18.66 7.86 ;
        RECT  14.94 4.14 15.42 7.86 ;
        RECT  14.94 4.14 15.96 4.62 ;
        RECT  15.48 3.00 15.96 4.62 ;
        RECT  15.90 5.10 16.50 5.70 ;
        RECT  14.88 8.34 15.48 8.94 ;
        RECT  13.50 3.00 14.94 3.48 ;
        RECT  13.74 6.18 14.34 6.78 ;
        RECT  13.80 4.02 14.28 6.78 ;
        RECT  13.74 4.02 14.34 4.62 ;
        RECT  11.46 9.54 11.94 12.36 ;
        RECT  11.70 4.14 12.18 10.02 ;
        RECT  11.58 7.26 12.18 7.86 ;
        RECT  11.58 7.32 13.20 7.80 ;
        RECT  11.46 3.00 11.94 4.62 ;
        RECT  5.82 7.38 6.30 12.36 ;
        RECT  5.82 8.46 10.20 8.94 ;
        RECT  9.72 7.38 10.20 8.94 ;
        RECT  9.72 7.38 11.10 7.86 ;
        RECT  5.70 3.00 6.18 7.86 ;
        RECT  8.82 2.94 9.42 3.54 ;
        RECT  7.26 4.02 7.86 4.62 ;
        RECT  7.26 7.26 7.86 7.86 ;
        RECT  6.66 2.94 7.26 3.54 ;
        RECT  4.80 10.68 5.28 12.36 ;
        RECT  4.74 11.58 5.34 12.18 ;
        RECT  4.62 2.94 5.22 3.54 ;
        RECT  3.60 9.54 4.08 12.36 ;
        RECT  3.60 9.54 4.62 10.02 ;
        RECT  4.14 4.14 4.62 10.02 ;
        RECT  4.02 6.18 4.62 6.78 ;
        RECT  3.54 4.14 4.62 4.62 ;
        RECT  3.54 3.00 4.02 4.62 ;
        RECT  3.00 8.34 3.60 8.94 ;
        RECT  1.86 4.02 2.46 4.62 ;
        RECT  1.32 2.94 1.92 3.54 ;
        RECT  1.38 10.68 1.86 12.36 ;
        RECT  1.32 11.58 1.92 12.18 ;
        LAYER via ;
        RECT  16.02 5.22 16.38 5.58 ;
        RECT  15.00 8.46 15.36 8.82 ;
        RECT  13.86 4.14 14.22 4.50 ;
        RECT  13.86 6.30 14.22 6.66 ;
        RECT  11.70 7.38 12.06 7.74 ;
        RECT  8.94 3.06 9.30 3.42 ;
        RECT  7.38 4.14 7.74 4.50 ;
        RECT  7.38 7.38 7.74 7.74 ;
        RECT  6.78 3.06 7.14 3.42 ;
        RECT  4.86 11.70 5.22 12.06 ;
        RECT  4.74 3.06 5.10 3.42 ;
        RECT  4.14 6.30 4.50 6.66 ;
        RECT  3.12 8.46 3.48 8.82 ;
        RECT  1.98 4.14 2.34 4.50 ;
        RECT  1.44 3.06 1.80 3.42 ;
        RECT  1.44 11.70 1.80 12.06 ;
        LAYER metal2 ;
        RECT  15.90 5.10 16.50 5.70 ;
        RECT  15.96 4.08 16.44 5.70 ;
        RECT  13.74 4.02 14.34 4.62 ;
        RECT  13.74 4.08 16.44 4.56 ;
        RECT  14.88 8.34 15.48 8.94 ;
        RECT  3.00 8.34 3.60 8.94 ;
        RECT  3.00 8.40 15.48 8.88 ;
        RECT  13.74 6.18 14.34 6.78 ;
        RECT  4.02 6.18 4.62 6.78 ;
        RECT  4.02 6.24 14.34 6.72 ;
        RECT  11.58 7.26 12.18 7.86 ;
        RECT  7.26 7.26 7.86 7.86 ;
        RECT  7.26 7.32 12.18 7.80 ;
        RECT  8.82 2.94 9.42 3.54 ;
        RECT  6.66 2.94 7.26 3.54 ;
        RECT  6.66 3.00 9.42 3.48 ;
        RECT  7.26 4.02 7.86 4.62 ;
        RECT  1.86 4.02 2.46 4.62 ;
        RECT  1.86 4.08 7.86 4.56 ;
        RECT  4.74 11.58 5.34 12.18 ;
        RECT  1.32 11.58 1.92 12.18 ;
        RECT  1.32 11.64 5.34 12.12 ;
        RECT  4.62 2.94 5.22 3.54 ;
        RECT  1.32 2.94 1.92 3.54 ;
        RECT  1.32 3.00 5.22 3.48 ;
    END
END dp_2

MACRO dp_4
    CLASS CORE ;
    FOREIGN dp_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.60 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  19.50 2.76 19.98 5.64 ;
        RECT  19.50 7.86 19.98 12.36 ;
        RECT  19.50 5.16 20.76 5.64 ;
        RECT  15.96 6.24 20.76 6.72 ;
        RECT  20.28 5.16 20.76 8.34 ;
        RECT  19.50 7.86 20.76 8.34 ;
        END
    END q
    PIN ip
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 7.32 1.32 7.80 ;
        END
    END ip
    PIN ck
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER metal1 ;
        RECT  3.00 6.24 3.48 6.72 ;
        END
    END ck
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.30 0.00 0.78 3.48 ;
        RECT  2.46 0.00 2.94 3.48 ;
        RECT  7.86 0.00 8.34 3.48 ;
        RECT  10.38 0.00 10.86 3.48 ;
        RECT  12.48 0.00 12.96 3.48 ;
        RECT  17.34 0.00 17.82 3.48 ;
        RECT  18.42 0.00 18.90 4.20 ;
        RECT  20.58 0.00 21.06 4.44 ;
        RECT  0.00 0.00 21.60 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.30 10.44 0.78 15.12 ;
        RECT  2.46 10.44 2.94 15.12 ;
        RECT  7.50 10.44 7.98 15.12 ;
        RECT  10.38 10.44 10.86 15.12 ;
        RECT  12.48 10.44 12.96 15.12 ;
        RECT  16.26 10.44 16.74 15.12 ;
        RECT  18.48 9.00 18.96 15.12 ;
        RECT  20.52 9.00 21.00 15.12 ;
        RECT  0.00 13.80 21.60 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  14.28 9.48 14.76 12.12 ;
        RECT  13.80 7.32 14.28 9.96 ;
        RECT  13.80 7.32 18.60 7.80 ;
        RECT  14.88 4.08 15.36 7.80 ;
        RECT  14.88 4.08 15.90 4.56 ;
        RECT  15.42 3.00 15.90 4.56 ;
        RECT  15.90 5.10 16.50 5.70 ;
        RECT  14.82 8.34 15.42 8.94 ;
        RECT  13.44 3.00 14.88 3.48 ;
        RECT  13.74 6.18 14.34 6.78 ;
        RECT  13.80 4.02 14.28 6.78 ;
        RECT  13.74 4.02 14.34 4.62 ;
        RECT  11.40 9.48 11.88 12.12 ;
        RECT  11.64 4.08 12.12 9.96 ;
        RECT  11.58 7.26 12.18 7.86 ;
        RECT  11.58 7.32 13.20 7.80 ;
        RECT  11.40 3.00 11.88 4.56 ;
        RECT  5.76 7.32 6.24 12.12 ;
        RECT  5.76 8.40 10.14 8.88 ;
        RECT  9.66 7.32 10.14 8.88 ;
        RECT  9.66 7.32 11.04 7.80 ;
        RECT  5.64 3.00 6.12 7.80 ;
        RECT  8.76 2.94 9.36 3.54 ;
        RECT  7.26 4.02 7.86 4.62 ;
        RECT  7.26 7.26 7.86 7.86 ;
        RECT  6.60 2.94 7.20 3.54 ;
        RECT  4.68 11.58 5.28 12.18 ;
        RECT  4.74 10.44 5.22 12.18 ;
        RECT  4.56 2.94 5.16 3.54 ;
        RECT  3.54 9.48 4.02 12.12 ;
        RECT  3.54 9.48 4.56 9.96 ;
        RECT  4.08 4.08 4.56 9.96 ;
        RECT  4.02 6.18 4.62 6.78 ;
        RECT  3.48 4.08 4.56 4.56 ;
        RECT  3.48 3.00 3.96 4.56 ;
        RECT  2.94 8.34 3.54 8.94 ;
        RECT  1.86 4.02 2.46 4.62 ;
        RECT  1.26 2.94 1.86 3.54 ;
        RECT  1.26 11.58 1.86 12.18 ;
        RECT  1.32 10.44 1.80 12.18 ;
        LAYER via ;
        RECT  16.02 5.22 16.38 5.58 ;
        RECT  14.94 8.46 15.30 8.82 ;
        RECT  13.86 4.14 14.22 4.50 ;
        RECT  13.86 6.30 14.22 6.66 ;
        RECT  11.70 7.38 12.06 7.74 ;
        RECT  8.88 3.06 9.24 3.42 ;
        RECT  7.38 4.14 7.74 4.50 ;
        RECT  7.38 7.38 7.74 7.74 ;
        RECT  6.72 3.06 7.08 3.42 ;
        RECT  4.80 11.70 5.16 12.06 ;
        RECT  4.68 3.06 5.04 3.42 ;
        RECT  4.14 6.30 4.50 6.66 ;
        RECT  3.06 8.46 3.42 8.82 ;
        RECT  1.98 4.14 2.34 4.50 ;
        RECT  1.38 3.06 1.74 3.42 ;
        RECT  1.38 11.70 1.74 12.06 ;
        LAYER metal2 ;
        RECT  15.90 5.10 16.50 5.70 ;
        RECT  15.96 4.08 16.44 5.70 ;
        RECT  13.74 4.02 14.34 4.62 ;
        RECT  13.74 4.08 16.44 4.56 ;
        RECT  14.82 8.34 15.42 8.94 ;
        RECT  2.94 8.34 3.54 8.94 ;
        RECT  2.94 8.40 15.42 8.88 ;
        RECT  13.74 6.18 14.34 6.78 ;
        RECT  4.02 6.18 4.62 6.78 ;
        RECT  4.02 6.24 14.34 6.72 ;
        RECT  11.58 7.26 12.18 7.86 ;
        RECT  7.26 7.26 7.86 7.86 ;
        RECT  7.26 7.32 12.18 7.80 ;
        RECT  8.76 2.94 9.36 3.54 ;
        RECT  6.60 2.94 7.20 3.54 ;
        RECT  6.60 3.00 9.36 3.48 ;
        RECT  7.26 4.02 7.86 4.62 ;
        RECT  1.86 4.02 2.46 4.62 ;
        RECT  1.86 4.08 7.86 4.56 ;
        RECT  4.68 11.58 5.28 12.18 ;
        RECT  1.26 11.58 1.86 12.18 ;
        RECT  1.26 11.64 5.28 12.12 ;
        RECT  4.56 2.94 5.16 3.54 ;
        RECT  1.26 2.94 1.86 3.54 ;
        RECT  1.26 3.00 5.16 3.48 ;
    END
END dp_4

MACRO drp_1
    CLASS CORE ;
    FOREIGN drp_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.76 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN rb
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal2 ;
        RECT  1.86 9.42 2.46 10.02 ;
        RECT  9.42 9.42 10.02 10.02 ;
        RECT  1.86 9.48 18.66 9.96 ;
        RECT  18.06 9.42 18.66 10.02 ;
        LAYER metal1 ;
        RECT  1.86 9.42 2.46 10.02 ;
        RECT  9.42 9.42 10.02 10.02 ;
        RECT  18.06 9.42 18.66 10.02 ;
        LAYER via ;
        RECT  1.98 9.54 2.34 9.90 ;
        RECT  9.54 9.54 9.90 9.90 ;
        RECT  18.18 9.54 18.54 9.90 ;
        END
    END rb
    PIN q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  21.36 6.24 22.92 6.72 ;
        RECT  22.44 4.08 22.92 12.12 ;
        RECT  22.56 3.00 23.04 4.56 ;
        END
    END q
    PIN ip
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 7.32 1.32 7.80 ;
        END
    END ip
    PIN ck
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER metal1 ;
        RECT  4.08 6.24 4.56 6.72 ;
        END
    END ck
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.60 0.00 1.08 3.48 ;
        RECT  3.54 0.00 4.02 3.48 ;
        RECT  8.94 0.00 9.42 3.48 ;
        RECT  12.54 0.00 13.02 3.48 ;
        RECT  14.64 0.00 15.12 3.48 ;
        RECT  21.42 0.00 21.90 3.48 ;
        RECT  0.00 0.00 23.76 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.30 10.44 0.78 15.12 ;
        RECT  2.28 10.44 2.76 15.12 ;
        RECT  3.36 10.44 3.84 15.12 ;
        RECT  8.88 10.44 9.36 15.12 ;
        RECT  12.54 10.44 13.02 15.12 ;
        RECT  14.64 10.44 15.12 15.12 ;
        RECT  18.60 10.44 19.08 15.12 ;
        RECT  21.36 10.44 21.84 15.12 ;
        RECT  0.00 13.80 23.76 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  16.44 9.48 16.92 12.12 ;
        RECT  15.96 7.32 16.44 9.96 ;
        RECT  15.96 7.32 21.84 7.80 ;
        RECT  17.04 4.08 17.52 7.80 ;
        RECT  17.04 4.08 18.06 4.56 ;
        RECT  17.58 3.00 18.06 4.56 ;
        RECT  19.38 3.00 20.88 3.48 ;
        RECT  20.28 11.58 20.88 12.18 ;
        RECT  20.34 10.44 20.82 12.18 ;
        RECT  18.06 5.10 18.66 5.70 ;
        RECT  17.52 11.58 18.12 12.18 ;
        RECT  17.58 10.44 18.06 12.18 ;
        RECT  16.98 8.34 17.58 8.94 ;
        RECT  15.60 3.00 17.04 3.48 ;
        RECT  15.90 6.18 16.50 6.78 ;
        RECT  15.96 4.02 16.44 6.78 ;
        RECT  15.90 4.02 16.50 4.62 ;
        RECT  13.56 9.48 14.04 12.12 ;
        RECT  13.80 4.08 14.28 9.96 ;
        RECT  13.74 7.26 14.34 7.86 ;
        RECT  13.74 7.32 15.36 7.80 ;
        RECT  13.56 3.00 14.04 4.56 ;
        RECT  6.84 7.32 7.32 12.12 ;
        RECT  6.84 8.40 12.30 8.88 ;
        RECT  11.82 7.32 12.30 8.88 ;
        RECT  11.82 7.32 13.20 7.80 ;
        RECT  6.72 3.00 7.20 7.80 ;
        RECT  10.92 2.94 11.52 3.54 ;
        RECT  9.90 11.58 10.50 12.18 ;
        RECT  9.96 10.44 10.44 12.18 ;
        RECT  8.34 4.02 8.94 4.62 ;
        RECT  8.34 7.26 8.94 7.86 ;
        RECT  7.80 11.58 8.40 12.18 ;
        RECT  7.86 10.44 8.34 12.18 ;
        RECT  7.68 2.94 8.28 3.54 ;
        RECT  5.76 11.58 6.36 12.18 ;
        RECT  5.82 10.44 6.30 12.18 ;
        RECT  5.64 2.94 6.24 3.54 ;
        RECT  4.44 9.48 4.92 12.12 ;
        RECT  4.44 9.48 5.64 9.96 ;
        RECT  5.16 4.08 5.64 9.96 ;
        RECT  5.10 6.18 5.70 6.78 ;
        RECT  4.56 4.08 5.64 4.56 ;
        RECT  4.56 3.00 5.04 4.56 ;
        RECT  4.02 8.34 4.62 8.94 ;
        RECT  2.94 4.02 3.54 4.62 ;
        RECT  2.28 2.94 2.88 3.54 ;
        RECT  1.26 11.58 1.86 12.18 ;
        RECT  1.32 10.44 1.80 12.18 ;
        LAYER via ;
        RECT  20.40 11.70 20.76 12.06 ;
        RECT  18.18 5.22 18.54 5.58 ;
        RECT  17.64 11.70 18.00 12.06 ;
        RECT  17.10 8.46 17.46 8.82 ;
        RECT  16.02 4.14 16.38 4.50 ;
        RECT  16.02 6.30 16.38 6.66 ;
        RECT  13.86 7.38 14.22 7.74 ;
        RECT  11.04 3.06 11.40 3.42 ;
        RECT  10.02 11.70 10.38 12.06 ;
        RECT  8.46 4.14 8.82 4.50 ;
        RECT  8.46 7.38 8.82 7.74 ;
        RECT  7.92 11.70 8.28 12.06 ;
        RECT  7.80 3.06 8.16 3.42 ;
        RECT  5.88 11.70 6.24 12.06 ;
        RECT  5.76 3.06 6.12 3.42 ;
        RECT  5.22 6.30 5.58 6.66 ;
        RECT  4.14 8.46 4.50 8.82 ;
        RECT  3.06 4.14 3.42 4.50 ;
        RECT  2.40 3.06 2.76 3.42 ;
        RECT  1.38 11.70 1.74 12.06 ;
        LAYER metal2 ;
        RECT  20.28 11.58 20.88 12.18 ;
        RECT  17.52 11.58 18.12 12.18 ;
        RECT  17.52 11.64 20.88 12.12 ;
        RECT  18.06 5.10 18.66 5.70 ;
        RECT  18.12 4.08 18.60 5.70 ;
        RECT  15.90 4.02 16.50 4.62 ;
        RECT  15.90 4.08 18.60 4.56 ;
        RECT  16.98 8.34 17.58 8.94 ;
        RECT  4.02 8.34 4.62 8.94 ;
        RECT  4.02 8.40 17.58 8.88 ;
        RECT  15.90 6.18 16.50 6.78 ;
        RECT  5.10 6.18 5.70 6.78 ;
        RECT  5.10 6.24 16.50 6.72 ;
        RECT  13.74 7.26 14.34 7.86 ;
        RECT  8.34 7.26 8.94 7.86 ;
        RECT  8.34 7.32 14.34 7.80 ;
        RECT  10.92 2.94 11.52 3.54 ;
        RECT  7.68 2.94 8.28 3.54 ;
        RECT  7.68 3.00 11.52 3.48 ;
        RECT  9.90 11.58 10.50 12.18 ;
        RECT  7.80 11.58 8.40 12.18 ;
        RECT  7.80 11.64 10.50 12.12 ;
        RECT  8.34 4.02 8.94 4.62 ;
        RECT  2.94 4.02 3.54 4.62 ;
        RECT  2.94 4.08 8.94 4.56 ;
        RECT  5.76 11.58 6.36 12.18 ;
        RECT  1.26 11.58 1.86 12.18 ;
        RECT  1.26 11.64 6.36 12.12 ;
        RECT  5.64 2.94 6.24 3.54 ;
        RECT  2.28 2.94 2.88 3.54 ;
        RECT  2.28 3.00 6.24 3.48 ;
    END
END drp_1

MACRO drp_2
    CLASS CORE ;
    FOREIGN drp_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.76 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN rb
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal2 ;
        RECT  1.86 9.42 2.46 10.02 ;
        RECT  9.42 9.42 10.02 10.02 ;
        RECT  1.86 9.48 18.66 9.96 ;
        RECT  18.06 9.42 18.66 10.02 ;
        LAYER metal1 ;
        RECT  1.86 9.42 2.46 10.02 ;
        RECT  9.42 9.42 10.02 10.02 ;
        RECT  18.06 9.42 18.66 10.02 ;
        LAYER via ;
        RECT  1.98 9.54 2.34 9.90 ;
        RECT  9.54 9.54 9.90 9.90 ;
        RECT  18.18 9.54 18.54 9.90 ;
        END
    END rb
    PIN q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  21.36 6.24 22.92 6.72 ;
        RECT  22.44 4.08 22.92 12.36 ;
        RECT  22.56 2.76 23.04 4.56 ;
        END
    END q
    PIN ip
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 7.32 1.32 7.80 ;
        END
    END ip
    PIN ck
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER metal1 ;
        RECT  4.08 6.24 4.56 6.72 ;
        END
    END ck
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.60 0.00 1.08 3.48 ;
        RECT  3.54 0.00 4.02 3.48 ;
        RECT  8.94 0.00 9.42 3.48 ;
        RECT  12.54 0.00 13.02 3.48 ;
        RECT  14.64 0.00 15.12 3.48 ;
        RECT  21.42 0.00 21.90 4.44 ;
        RECT  0.00 0.00 23.76 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.30 10.44 0.78 15.12 ;
        RECT  2.28 10.44 2.76 15.12 ;
        RECT  3.36 10.44 3.84 15.12 ;
        RECT  8.88 10.44 9.36 15.12 ;
        RECT  12.54 10.44 13.02 15.12 ;
        RECT  14.64 10.44 15.12 15.12 ;
        RECT  18.60 10.44 19.08 15.12 ;
        RECT  21.36 9.00 21.84 15.12 ;
        RECT  0.00 13.80 23.76 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  16.44 9.48 16.92 12.12 ;
        RECT  15.96 7.32 16.44 9.96 ;
        RECT  15.96 7.32 21.84 7.80 ;
        RECT  17.04 4.08 17.52 7.80 ;
        RECT  17.04 4.08 18.06 4.56 ;
        RECT  17.58 3.00 18.06 4.56 ;
        RECT  20.40 2.76 20.88 4.44 ;
        RECT  19.38 3.00 20.88 3.48 ;
        RECT  20.28 11.58 20.88 12.18 ;
        RECT  20.34 9.00 20.82 12.18 ;
        RECT  18.06 5.10 18.66 5.70 ;
        RECT  17.52 11.58 18.12 12.18 ;
        RECT  17.58 10.44 18.06 12.18 ;
        RECT  16.98 8.34 17.58 8.94 ;
        RECT  15.60 3.00 17.04 3.48 ;
        RECT  15.90 6.18 16.50 6.78 ;
        RECT  15.96 4.02 16.44 6.78 ;
        RECT  15.90 4.02 16.50 4.62 ;
        RECT  13.56 9.48 14.04 12.12 ;
        RECT  13.80 4.08 14.28 9.96 ;
        RECT  13.74 7.26 14.34 7.86 ;
        RECT  13.74 7.32 15.36 7.80 ;
        RECT  13.56 3.00 14.04 4.56 ;
        RECT  6.84 7.32 7.32 12.12 ;
        RECT  6.84 8.40 12.30 8.88 ;
        RECT  11.82 7.32 12.30 8.88 ;
        RECT  11.82 7.32 13.20 7.80 ;
        RECT  6.72 3.00 7.20 7.80 ;
        RECT  10.92 2.94 11.52 3.54 ;
        RECT  9.90 11.58 10.50 12.18 ;
        RECT  9.96 10.44 10.44 12.18 ;
        RECT  8.34 4.02 8.94 4.62 ;
        RECT  8.34 7.26 8.94 7.86 ;
        RECT  7.80 11.58 8.40 12.18 ;
        RECT  7.86 10.44 8.34 12.18 ;
        RECT  7.68 2.94 8.28 3.54 ;
        RECT  5.76 11.52 6.36 12.12 ;
        RECT  5.82 10.44 6.30 12.12 ;
        RECT  5.64 2.94 6.24 3.54 ;
        RECT  4.44 9.48 4.92 12.12 ;
        RECT  4.44 9.48 5.64 9.96 ;
        RECT  5.16 4.08 5.64 9.96 ;
        RECT  5.10 6.18 5.70 6.78 ;
        RECT  4.56 4.08 5.64 4.56 ;
        RECT  4.56 3.00 5.04 4.56 ;
        RECT  4.02 8.34 4.62 8.94 ;
        RECT  2.94 4.02 3.54 4.62 ;
        RECT  2.28 2.94 2.88 3.54 ;
        RECT  1.26 11.58 1.86 12.18 ;
        RECT  1.32 10.44 1.80 12.18 ;
        LAYER via ;
        RECT  20.40 11.70 20.76 12.06 ;
        RECT  18.18 5.22 18.54 5.58 ;
        RECT  17.64 11.70 18.00 12.06 ;
        RECT  17.10 8.46 17.46 8.82 ;
        RECT  16.02 4.14 16.38 4.50 ;
        RECT  16.02 6.30 16.38 6.66 ;
        RECT  13.86 7.38 14.22 7.74 ;
        RECT  11.04 3.06 11.40 3.42 ;
        RECT  10.02 11.70 10.38 12.06 ;
        RECT  8.46 4.14 8.82 4.50 ;
        RECT  8.46 7.38 8.82 7.74 ;
        RECT  7.92 11.70 8.28 12.06 ;
        RECT  7.80 3.06 8.16 3.42 ;
        RECT  5.88 11.64 6.24 12.00 ;
        RECT  5.76 3.06 6.12 3.42 ;
        RECT  5.22 6.30 5.58 6.66 ;
        RECT  4.14 8.46 4.50 8.82 ;
        RECT  3.06 4.14 3.42 4.50 ;
        RECT  2.40 3.06 2.76 3.42 ;
        RECT  1.38 11.70 1.74 12.06 ;
        LAYER metal2 ;
        RECT  20.28 11.58 20.88 12.18 ;
        RECT  17.52 11.58 18.12 12.18 ;
        RECT  17.52 11.64 20.88 12.12 ;
        RECT  18.06 5.10 18.66 5.70 ;
        RECT  18.12 4.08 18.60 5.70 ;
        RECT  15.90 4.02 16.50 4.62 ;
        RECT  15.90 4.08 18.60 4.56 ;
        RECT  16.98 8.34 17.58 8.94 ;
        RECT  4.02 8.34 4.62 8.94 ;
        RECT  4.02 8.40 17.58 8.88 ;
        RECT  15.90 6.18 16.50 6.78 ;
        RECT  5.10 6.18 5.70 6.78 ;
        RECT  5.10 6.24 16.50 6.72 ;
        RECT  13.74 7.26 14.34 7.86 ;
        RECT  8.34 7.26 8.94 7.86 ;
        RECT  8.34 7.32 14.34 7.80 ;
        RECT  10.92 2.94 11.52 3.54 ;
        RECT  7.68 2.94 8.28 3.54 ;
        RECT  7.68 3.00 11.52 3.48 ;
        RECT  9.90 11.58 10.50 12.18 ;
        RECT  7.80 11.58 8.40 12.18 ;
        RECT  7.80 11.64 10.50 12.12 ;
        RECT  8.34 4.02 8.94 4.62 ;
        RECT  2.94 4.02 3.54 4.62 ;
        RECT  2.94 4.08 8.94 4.56 ;
        RECT  1.26 11.58 1.86 12.18 ;
        RECT  1.26 11.64 6.36 12.12 ;
        RECT  5.76 11.52 6.36 12.12 ;
        RECT  5.64 2.94 6.24 3.54 ;
        RECT  2.28 2.94 2.88 3.54 ;
        RECT  2.28 3.00 6.24 3.48 ;
    END
END drp_2

MACRO drp_4
    CLASS CORE ;
    FOREIGN drp_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 24.84 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN rb
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal2 ;
        RECT  1.86 9.42 2.46 10.02 ;
        RECT  9.42 9.42 10.02 10.02 ;
        RECT  1.86 9.48 18.66 9.96 ;
        RECT  18.06 9.42 18.66 10.02 ;
        LAYER metal1 ;
        RECT  1.86 9.42 2.46 10.02 ;
        RECT  9.42 9.42 10.02 10.02 ;
        RECT  18.06 9.42 18.66 10.02 ;
        LAYER via ;
        RECT  1.98 9.54 2.34 9.90 ;
        RECT  9.54 9.54 9.90 9.90 ;
        RECT  18.18 9.54 18.54 9.90 ;
        END
    END rb
    PIN q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  21.36 6.24 22.92 6.72 ;
        RECT  22.44 4.08 22.92 12.36 ;
        RECT  22.50 2.76 22.98 4.56 ;
        END
    END q
    PIN ip
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 7.32 1.32 7.80 ;
        END
    END ip
    PIN ck
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER metal1 ;
        RECT  4.08 6.24 4.56 6.72 ;
        END
    END ck
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.60 0.00 1.08 3.48 ;
        RECT  3.54 0.00 4.02 3.48 ;
        RECT  8.94 0.00 9.42 3.48 ;
        RECT  12.54 0.00 13.02 3.48 ;
        RECT  14.64 0.00 15.12 3.48 ;
        RECT  21.42 0.00 21.90 4.44 ;
        RECT  23.64 0.00 24.12 4.44 ;
        RECT  0.00 0.00 24.84 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.30 10.44 0.78 15.12 ;
        RECT  2.28 10.44 2.76 15.12 ;
        RECT  3.36 10.44 3.84 15.12 ;
        RECT  8.88 10.44 9.36 15.12 ;
        RECT  12.54 10.44 13.02 15.12 ;
        RECT  14.64 10.44 15.12 15.12 ;
        RECT  18.60 10.44 19.08 15.12 ;
        RECT  21.36 9.00 21.84 15.12 ;
        RECT  23.58 9.00 24.06 15.12 ;
        RECT  0.00 13.80 24.84 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  16.44 9.48 16.92 12.12 ;
        RECT  15.96 7.32 16.44 9.96 ;
        RECT  15.96 7.32 21.84 7.80 ;
        RECT  17.04 4.08 17.52 7.80 ;
        RECT  17.04 4.08 18.06 4.56 ;
        RECT  17.58 3.00 18.06 4.56 ;
        RECT  20.40 2.76 20.88 4.44 ;
        RECT  19.38 3.00 20.88 3.48 ;
        RECT  20.28 11.58 20.88 12.18 ;
        RECT  20.34 9.00 20.82 12.18 ;
        RECT  18.06 5.10 18.66 5.70 ;
        RECT  17.52 11.58 18.12 12.18 ;
        RECT  17.58 10.44 18.06 12.18 ;
        RECT  16.98 8.34 17.58 8.94 ;
        RECT  15.60 3.00 17.04 3.48 ;
        RECT  15.90 6.18 16.50 6.78 ;
        RECT  15.96 4.02 16.44 6.78 ;
        RECT  15.90 4.02 16.50 4.62 ;
        RECT  13.56 9.48 14.04 12.12 ;
        RECT  13.80 4.08 14.28 9.96 ;
        RECT  13.74 7.26 14.34 7.86 ;
        RECT  13.74 7.32 15.36 7.80 ;
        RECT  13.56 3.00 14.04 4.56 ;
        RECT  6.84 7.32 7.32 12.12 ;
        RECT  6.84 8.40 12.30 8.88 ;
        RECT  11.82 7.32 12.30 8.88 ;
        RECT  11.82 7.32 13.20 7.80 ;
        RECT  6.72 3.00 7.20 7.80 ;
        RECT  10.92 2.94 11.52 3.54 ;
        RECT  9.90 11.58 10.50 12.18 ;
        RECT  9.96 10.44 10.44 12.18 ;
        RECT  8.34 4.02 8.94 4.62 ;
        RECT  8.34 7.26 8.94 7.86 ;
        RECT  7.80 11.58 8.40 12.18 ;
        RECT  7.86 10.44 8.34 12.18 ;
        RECT  7.68 2.94 8.28 3.54 ;
        RECT  5.76 11.58 6.36 12.18 ;
        RECT  5.82 10.44 6.30 12.18 ;
        RECT  5.64 2.94 6.24 3.54 ;
        RECT  4.44 9.48 4.92 12.12 ;
        RECT  4.44 9.48 5.64 9.96 ;
        RECT  5.16 4.08 5.64 9.96 ;
        RECT  5.10 6.18 5.70 6.78 ;
        RECT  4.56 4.08 5.64 4.56 ;
        RECT  4.56 3.00 5.04 4.56 ;
        RECT  4.02 8.34 4.62 8.94 ;
        RECT  2.94 4.02 3.54 4.62 ;
        RECT  2.28 2.94 2.88 3.54 ;
        RECT  1.26 11.58 1.86 12.18 ;
        RECT  1.32 10.44 1.80 12.18 ;
        LAYER via ;
        RECT  20.40 11.70 20.76 12.06 ;
        RECT  18.18 5.22 18.54 5.58 ;
        RECT  17.64 11.70 18.00 12.06 ;
        RECT  17.10 8.46 17.46 8.82 ;
        RECT  16.02 4.14 16.38 4.50 ;
        RECT  16.02 6.30 16.38 6.66 ;
        RECT  13.86 7.38 14.22 7.74 ;
        RECT  11.04 3.06 11.40 3.42 ;
        RECT  10.02 11.70 10.38 12.06 ;
        RECT  8.46 4.14 8.82 4.50 ;
        RECT  8.46 7.38 8.82 7.74 ;
        RECT  7.92 11.70 8.28 12.06 ;
        RECT  7.80 3.06 8.16 3.42 ;
        RECT  5.88 11.70 6.24 12.06 ;
        RECT  5.76 3.06 6.12 3.42 ;
        RECT  5.22 6.30 5.58 6.66 ;
        RECT  4.14 8.46 4.50 8.82 ;
        RECT  3.06 4.14 3.42 4.50 ;
        RECT  2.40 3.06 2.76 3.42 ;
        RECT  1.38 11.70 1.74 12.06 ;
        LAYER metal2 ;
        RECT  20.28 11.58 20.88 12.18 ;
        RECT  17.52 11.58 18.12 12.18 ;
        RECT  17.52 11.64 20.88 12.12 ;
        RECT  18.06 5.10 18.66 5.70 ;
        RECT  18.12 4.08 18.60 5.70 ;
        RECT  15.90 4.02 16.50 4.62 ;
        RECT  15.90 4.08 18.60 4.56 ;
        RECT  16.98 8.34 17.58 8.94 ;
        RECT  4.02 8.34 4.62 8.94 ;
        RECT  4.02 8.40 17.58 8.88 ;
        RECT  15.90 6.18 16.50 6.78 ;
        RECT  5.10 6.18 5.70 6.78 ;
        RECT  5.10 6.18 16.50 6.66 ;
        RECT  13.74 7.26 14.34 7.86 ;
        RECT  8.34 7.26 8.94 7.86 ;
        RECT  8.34 7.32 14.34 7.80 ;
        RECT  10.92 2.94 11.52 3.54 ;
        RECT  7.68 2.94 8.28 3.54 ;
        RECT  7.68 3.00 11.52 3.48 ;
        RECT  9.90 11.58 10.50 12.18 ;
        RECT  7.80 11.58 8.40 12.18 ;
        RECT  7.80 11.64 10.50 12.12 ;
        RECT  8.34 4.02 8.94 4.62 ;
        RECT  2.94 4.02 3.54 4.62 ;
        RECT  2.94 4.08 8.94 4.56 ;
        RECT  5.76 11.58 6.36 12.18 ;
        RECT  1.26 11.58 1.86 12.18 ;
        RECT  1.26 11.64 6.36 12.12 ;
        RECT  5.64 2.94 6.24 3.54 ;
        RECT  2.28 2.94 2.88 3.54 ;
        RECT  2.28 3.00 6.24 3.48 ;
    END
END drp_4

MACRO drsp_1
    CLASS CORE ;
    FOREIGN drsp_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 27.00 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN s
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal2 ;
        RECT  1.86 5.10 2.46 5.70 ;
        RECT  9.42 5.10 10.02 5.70 ;
        RECT  1.86 5.16 19.68 5.64 ;
        RECT  19.20 5.16 19.68 6.72 ;
        RECT  19.20 6.24 22.98 6.72 ;
        RECT  22.38 6.18 22.98 6.78 ;
        LAYER metal1 ;
        RECT  1.86 5.10 2.46 5.70 ;
        RECT  9.42 5.10 10.02 5.70 ;
        RECT  22.38 6.18 22.98 6.78 ;
        LAYER via ;
        RECT  1.98 5.22 2.34 5.58 ;
        RECT  9.54 5.22 9.90 5.58 ;
        RECT  22.50 6.30 22.86 6.66 ;
        END
    END s
    PIN rb
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal2 ;
        RECT  2.94 9.42 3.54 10.02 ;
        RECT  11.58 9.42 12.18 10.02 ;
        RECT  2.94 9.48 20.82 9.96 ;
        RECT  20.22 9.42 20.82 10.02 ;
        LAYER metal1 ;
        RECT  2.94 9.42 3.54 10.02 ;
        RECT  11.58 9.42 12.18 10.02 ;
        RECT  20.22 9.42 20.82 10.02 ;
        LAYER via ;
        RECT  3.06 9.54 3.42 9.90 ;
        RECT  11.70 9.54 12.06 9.90 ;
        RECT  20.34 9.54 20.70 9.90 ;
        END
    END rb
    PIN q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  24.60 6.24 26.16 6.72 ;
        RECT  25.32 9.48 25.80 12.12 ;
        RECT  25.56 3.00 26.04 4.56 ;
        RECT  25.68 4.08 26.16 9.96 ;
        END
    END q
    PIN ip
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 7.32 1.32 7.80 ;
        END
    END ip
    PIN ck
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER metal1 ;
        RECT  5.16 6.24 5.64 6.72 ;
        END
    END ck
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.38 0.00 1.86 3.48 ;
        RECT  4.62 0.00 5.10 3.48 ;
        RECT  11.52 0.00 12.00 3.48 ;
        RECT  14.70 0.00 15.18 3.48 ;
        RECT  16.80 0.00 17.28 3.48 ;
        RECT  22.50 0.00 22.98 3.48 ;
        RECT  24.54 0.00 25.02 3.48 ;
        RECT  0.00 0.00 27.00 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.66 10.44 1.14 15.12 ;
        RECT  3.36 10.44 3.84 15.12 ;
        RECT  4.44 10.44 4.92 15.12 ;
        RECT  10.80 10.44 11.28 15.12 ;
        RECT  14.70 10.44 15.18 15.12 ;
        RECT  16.80 10.44 17.28 15.12 ;
        RECT  20.76 10.44 21.24 15.12 ;
        RECT  24.24 10.44 24.72 15.12 ;
        RECT  0.00 13.80 27.00 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  18.60 9.48 19.08 12.12 ;
        RECT  18.12 7.32 18.60 9.96 ;
        RECT  18.12 7.32 25.08 7.80 ;
        RECT  19.20 4.08 19.68 7.80 ;
        RECT  19.20 4.08 20.22 4.56 ;
        RECT  19.74 3.00 20.22 4.56 ;
        RECT  21.54 4.20 24.06 4.68 ;
        RECT  23.58 3.00 24.06 4.68 ;
        RECT  21.54 3.00 22.02 4.68 ;
        RECT  22.38 11.58 22.98 12.18 ;
        RECT  22.50 10.44 22.98 12.18 ;
        RECT  20.22 5.10 20.82 5.70 ;
        RECT  19.68 11.58 20.28 12.18 ;
        RECT  19.74 10.44 20.22 12.18 ;
        RECT  19.14 8.34 19.74 8.94 ;
        RECT  17.76 3.00 19.20 3.48 ;
        RECT  18.06 6.18 18.66 6.78 ;
        RECT  18.12 4.02 18.60 6.78 ;
        RECT  18.06 4.02 18.66 4.62 ;
        RECT  15.72 9.48 16.20 12.12 ;
        RECT  15.96 4.08 16.44 9.96 ;
        RECT  15.90 7.26 16.50 7.86 ;
        RECT  15.90 7.32 17.52 7.80 ;
        RECT  15.72 3.00 16.20 4.56 ;
        RECT  7.92 7.32 8.40 12.12 ;
        RECT  7.92 8.40 14.46 8.88 ;
        RECT  13.98 7.32 14.46 8.88 ;
        RECT  13.98 7.32 15.36 7.80 ;
        RECT  7.80 3.00 8.28 7.80 ;
        RECT  13.50 2.94 14.10 3.54 ;
        RECT  10.56 4.08 12.96 4.56 ;
        RECT  12.48 3.00 12.96 4.56 ;
        RECT  10.56 3.00 11.04 4.56 ;
        RECT  11.76 11.58 12.36 12.18 ;
        RECT  11.82 10.44 12.30 12.18 ;
        RECT  10.50 7.26 11.10 7.86 ;
        RECT  9.42 4.02 10.02 4.62 ;
        RECT  8.88 11.58 9.48 12.18 ;
        RECT  8.94 10.44 9.42 12.18 ;
        RECT  8.76 2.94 9.36 3.54 ;
        RECT  6.84 11.58 7.44 12.18 ;
        RECT  6.90 10.44 7.38 12.18 ;
        RECT  6.72 2.94 7.32 3.54 ;
        RECT  5.52 9.48 6.00 12.12 ;
        RECT  5.52 9.48 6.72 9.96 ;
        RECT  6.24 4.08 6.72 9.96 ;
        RECT  6.18 6.18 6.78 6.78 ;
        RECT  5.64 4.08 6.72 4.56 ;
        RECT  5.64 3.00 6.12 4.56 ;
        RECT  5.10 8.34 5.70 8.94 ;
        RECT  4.02 4.02 4.62 4.62 ;
        RECT  3.36 2.94 3.96 3.54 ;
        RECT  2.34 11.58 2.94 12.18 ;
        RECT  2.40 10.44 2.88 12.18 ;
        RECT  0.42 4.08 2.82 4.56 ;
        RECT  2.34 3.00 2.82 4.56 ;
        RECT  0.42 3.00 0.90 4.56 ;
        LAYER via ;
        RECT  22.50 11.70 22.86 12.06 ;
        RECT  20.34 5.22 20.70 5.58 ;
        RECT  19.80 11.70 20.16 12.06 ;
        RECT  19.26 8.46 19.62 8.82 ;
        RECT  18.18 4.14 18.54 4.50 ;
        RECT  18.18 6.30 18.54 6.66 ;
        RECT  16.02 7.38 16.38 7.74 ;
        RECT  13.62 3.06 13.98 3.42 ;
        RECT  11.88 11.70 12.24 12.06 ;
        RECT  10.62 7.38 10.98 7.74 ;
        RECT  9.54 4.14 9.90 4.50 ;
        RECT  9.00 11.70 9.36 12.06 ;
        RECT  8.88 3.06 9.24 3.42 ;
        RECT  6.96 11.70 7.32 12.06 ;
        RECT  6.84 3.06 7.20 3.42 ;
        RECT  6.30 6.30 6.66 6.66 ;
        RECT  5.22 8.46 5.58 8.82 ;
        RECT  4.14 4.14 4.50 4.50 ;
        RECT  3.48 3.06 3.84 3.42 ;
        RECT  2.46 11.70 2.82 12.06 ;
        LAYER metal2 ;
        RECT  22.38 11.58 22.98 12.18 ;
        RECT  19.68 11.58 20.28 12.18 ;
        RECT  19.68 11.64 22.98 12.12 ;
        RECT  20.22 5.10 20.82 5.70 ;
        RECT  20.28 4.08 20.76 5.70 ;
        RECT  18.06 4.02 18.66 4.62 ;
        RECT  18.06 4.08 20.76 4.56 ;
        RECT  19.14 8.34 19.74 8.94 ;
        RECT  5.10 8.34 5.70 8.94 ;
        RECT  5.10 8.40 19.74 8.88 ;
        RECT  18.06 6.18 18.66 6.78 ;
        RECT  6.18 6.18 6.78 6.78 ;
        RECT  6.18 6.24 18.66 6.72 ;
        RECT  15.90 7.26 16.50 7.86 ;
        RECT  10.50 7.26 11.10 7.86 ;
        RECT  10.50 7.32 16.50 7.80 ;
        RECT  13.50 2.94 14.10 3.54 ;
        RECT  8.76 2.94 9.36 3.54 ;
        RECT  8.76 3.00 14.10 3.48 ;
        RECT  11.76 11.58 12.36 12.18 ;
        RECT  8.88 11.58 9.48 12.18 ;
        RECT  8.88 11.64 12.36 12.12 ;
        RECT  9.42 4.02 10.02 4.62 ;
        RECT  4.02 4.02 4.62 4.62 ;
        RECT  4.02 4.08 10.02 4.56 ;
        RECT  6.84 11.58 7.44 12.18 ;
        RECT  2.34 11.58 2.94 12.18 ;
        RECT  2.34 11.64 7.44 12.12 ;
        RECT  6.72 2.94 7.32 3.54 ;
        RECT  3.36 2.94 3.96 3.54 ;
        RECT  3.36 3.00 7.32 3.48 ;
    END
END drsp_1

MACRO drsp_2
    CLASS CORE ;
    FOREIGN drsp_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 27.00 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN s
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal2 ;
        RECT  1.86 5.10 2.46 5.70 ;
        RECT  9.42 5.10 10.02 5.70 ;
        RECT  1.86 5.16 19.68 5.64 ;
        RECT  19.20 5.16 19.68 6.72 ;
        RECT  19.20 6.24 22.98 6.72 ;
        RECT  22.38 6.18 22.98 6.78 ;
        LAYER metal1 ;
        RECT  1.86 5.10 2.46 5.70 ;
        RECT  9.42 5.10 10.02 5.70 ;
        RECT  22.38 6.18 22.98 6.78 ;
        LAYER via ;
        RECT  1.98 5.22 2.34 5.58 ;
        RECT  9.54 5.22 9.90 5.58 ;
        RECT  22.50 6.30 22.86 6.66 ;
        END
    END s
    PIN rb
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal2 ;
        RECT  2.94 9.42 3.54 10.02 ;
        RECT  11.58 9.42 12.18 10.02 ;
        RECT  2.94 9.48 20.82 9.96 ;
        RECT  20.22 9.42 20.82 10.02 ;
        LAYER metal1 ;
        RECT  2.94 9.42 3.54 10.02 ;
        RECT  11.58 9.42 12.18 10.02 ;
        RECT  20.22 9.42 20.82 10.02 ;
        LAYER via ;
        RECT  3.06 9.54 3.42 9.90 ;
        RECT  11.70 9.54 12.06 9.90 ;
        RECT  20.34 9.54 20.70 9.90 ;
        END
    END rb
    PIN q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  24.60 6.24 26.16 6.72 ;
        RECT  25.32 8.40 25.80 12.36 ;
        RECT  25.56 2.76 26.04 4.56 ;
        RECT  25.68 4.08 26.16 8.88 ;
        END
    END q
    PIN ip
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 7.32 1.32 7.80 ;
        END
    END ip
    PIN ck
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER metal1 ;
        RECT  5.16 6.24 5.64 6.72 ;
        END
    END ck
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.38 0.00 1.86 3.48 ;
        RECT  4.62 0.00 5.10 3.48 ;
        RECT  11.52 0.00 12.00 3.48 ;
        RECT  14.70 0.00 15.18 3.48 ;
        RECT  16.80 0.00 17.28 3.48 ;
        RECT  22.50 0.00 22.98 4.44 ;
        RECT  24.54 0.00 25.02 4.44 ;
        RECT  0.00 0.00 27.00 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.66 10.44 1.14 15.12 ;
        RECT  3.36 10.44 3.84 15.12 ;
        RECT  4.44 10.44 4.92 15.12 ;
        RECT  10.80 10.44 11.28 15.12 ;
        RECT  14.70 10.44 15.18 15.12 ;
        RECT  16.80 10.44 17.28 15.12 ;
        RECT  20.76 10.44 21.24 15.12 ;
        RECT  24.24 9.00 24.72 15.12 ;
        RECT  0.00 13.80 27.00 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  18.60 9.48 19.08 12.12 ;
        RECT  18.12 7.32 18.60 9.96 ;
        RECT  18.12 7.32 25.08 7.80 ;
        RECT  19.20 4.08 19.68 7.80 ;
        RECT  19.20 4.08 20.22 4.56 ;
        RECT  19.74 3.00 20.22 4.56 ;
        RECT  21.54 5.16 24.06 5.64 ;
        RECT  23.58 2.76 24.06 5.64 ;
        RECT  21.54 3.00 22.02 5.64 ;
        RECT  22.50 9.00 22.98 12.36 ;
        RECT  22.38 11.58 22.98 12.18 ;
        RECT  20.22 5.10 20.82 5.70 ;
        RECT  19.68 11.58 20.28 12.18 ;
        RECT  19.74 10.44 20.22 12.18 ;
        RECT  19.14 8.34 19.74 8.94 ;
        RECT  17.76 3.00 19.20 3.48 ;
        RECT  18.06 6.18 18.66 6.78 ;
        RECT  18.12 4.02 18.60 6.78 ;
        RECT  18.06 4.02 18.66 4.62 ;
        RECT  15.72 9.48 16.20 12.12 ;
        RECT  15.96 4.08 16.44 9.96 ;
        RECT  15.90 7.26 16.50 7.86 ;
        RECT  15.90 7.32 17.52 7.80 ;
        RECT  15.72 3.00 16.20 4.56 ;
        RECT  7.92 7.32 8.40 12.36 ;
        RECT  7.92 8.40 14.46 8.88 ;
        RECT  13.98 7.32 14.46 8.88 ;
        RECT  13.98 7.32 15.36 7.80 ;
        RECT  7.80 3.00 8.28 7.80 ;
        RECT  13.50 2.94 14.10 3.54 ;
        RECT  10.56 4.08 12.96 4.56 ;
        RECT  12.48 3.00 12.96 4.56 ;
        RECT  10.56 3.00 11.04 4.56 ;
        RECT  11.76 11.58 12.36 12.18 ;
        RECT  11.82 10.44 12.30 12.18 ;
        RECT  10.50 7.26 11.10 7.86 ;
        RECT  9.42 4.02 10.02 4.62 ;
        RECT  8.88 11.58 9.48 12.18 ;
        RECT  8.94 10.44 9.42 12.18 ;
        RECT  8.76 2.94 9.36 3.54 ;
        RECT  6.84 11.58 7.44 12.18 ;
        RECT  6.90 10.44 7.38 12.18 ;
        RECT  6.72 2.94 7.32 3.54 ;
        RECT  5.52 9.48 6.00 12.12 ;
        RECT  5.52 9.48 6.72 9.96 ;
        RECT  6.24 4.08 6.72 9.96 ;
        RECT  6.18 6.18 6.78 6.78 ;
        RECT  5.64 4.08 6.72 4.56 ;
        RECT  5.64 3.00 6.12 4.56 ;
        RECT  5.10 8.34 5.70 8.94 ;
        RECT  4.02 4.02 4.62 4.62 ;
        RECT  3.36 2.94 3.96 3.54 ;
        RECT  2.34 11.58 2.94 12.18 ;
        RECT  2.40 10.44 2.88 12.18 ;
        RECT  0.42 4.08 2.82 4.56 ;
        RECT  2.34 3.00 2.82 4.56 ;
        RECT  0.42 3.00 0.90 4.56 ;
        LAYER via ;
        RECT  22.50 11.70 22.86 12.06 ;
        RECT  20.34 5.22 20.70 5.58 ;
        RECT  19.80 11.70 20.16 12.06 ;
        RECT  19.26 8.46 19.62 8.82 ;
        RECT  18.18 4.14 18.54 4.50 ;
        RECT  18.18 6.30 18.54 6.66 ;
        RECT  16.02 7.38 16.38 7.74 ;
        RECT  13.62 3.06 13.98 3.42 ;
        RECT  11.88 11.70 12.24 12.06 ;
        RECT  10.62 7.38 10.98 7.74 ;
        RECT  9.54 4.14 9.90 4.50 ;
        RECT  9.00 11.70 9.36 12.06 ;
        RECT  8.88 3.06 9.24 3.42 ;
        RECT  6.96 11.70 7.32 12.06 ;
        RECT  6.84 3.06 7.20 3.42 ;
        RECT  6.30 6.30 6.66 6.66 ;
        RECT  5.22 8.46 5.58 8.82 ;
        RECT  4.14 4.14 4.50 4.50 ;
        RECT  3.48 3.06 3.84 3.42 ;
        RECT  2.46 11.70 2.82 12.06 ;
        LAYER metal2 ;
        RECT  22.38 11.58 22.98 12.18 ;
        RECT  19.68 11.58 20.28 12.18 ;
        RECT  19.68 11.64 22.98 12.12 ;
        RECT  20.22 5.10 20.82 5.70 ;
        RECT  20.28 4.08 20.76 5.70 ;
        RECT  18.06 4.02 18.66 4.62 ;
        RECT  18.06 4.08 20.76 4.56 ;
        RECT  19.14 8.34 19.74 8.94 ;
        RECT  5.10 8.34 5.70 8.94 ;
        RECT  5.10 8.40 19.74 8.88 ;
        RECT  18.06 6.18 18.66 6.78 ;
        RECT  6.18 6.18 6.78 6.78 ;
        RECT  6.18 6.24 18.66 6.72 ;
        RECT  15.90 7.26 16.50 7.86 ;
        RECT  10.50 7.26 11.10 7.86 ;
        RECT  10.50 7.32 16.50 7.80 ;
        RECT  13.50 2.94 14.10 3.54 ;
        RECT  8.76 2.94 9.36 3.54 ;
        RECT  8.76 3.00 14.10 3.48 ;
        RECT  11.76 11.58 12.36 12.18 ;
        RECT  8.88 11.58 9.48 12.18 ;
        RECT  8.88 11.64 12.36 12.12 ;
        RECT  9.42 4.02 10.02 4.62 ;
        RECT  4.02 4.02 4.62 4.62 ;
        RECT  4.02 4.08 10.02 4.56 ;
        RECT  6.84 11.58 7.44 12.18 ;
        RECT  2.34 11.58 2.94 12.18 ;
        RECT  2.34 11.64 7.44 12.12 ;
        RECT  6.72 2.94 7.32 3.54 ;
        RECT  3.36 2.94 3.96 3.54 ;
        RECT  3.36 3.00 7.32 3.48 ;
    END
END drsp_2

MACRO drsp_4
    CLASS CORE ;
    FOREIGN drsp_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 28.08 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN s
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal2 ;
        RECT  1.86 5.10 2.46 5.70 ;
        RECT  9.42 5.10 10.02 5.70 ;
        RECT  1.86 5.16 19.68 5.64 ;
        RECT  19.20 5.16 19.68 6.72 ;
        RECT  19.20 6.24 22.98 6.72 ;
        RECT  22.38 6.18 22.98 6.78 ;
        LAYER metal1 ;
        RECT  1.86 5.10 2.46 5.70 ;
        RECT  9.42 5.10 10.02 5.70 ;
        RECT  22.38 6.18 22.98 6.78 ;
        LAYER via ;
        RECT  1.98 5.22 2.34 5.58 ;
        RECT  9.54 5.22 9.90 5.58 ;
        RECT  22.50 6.30 22.86 6.66 ;
        END
    END s
    PIN rb
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal2 ;
        RECT  2.94 9.42 3.54 10.02 ;
        RECT  11.58 9.42 12.18 10.02 ;
        RECT  2.94 9.48 20.82 9.96 ;
        RECT  20.22 9.42 20.82 10.02 ;
        LAYER metal1 ;
        RECT  2.94 9.42 3.54 10.02 ;
        RECT  11.58 9.42 12.18 10.02 ;
        RECT  20.22 9.42 20.82 10.02 ;
        LAYER via ;
        RECT  3.06 9.54 3.42 9.90 ;
        RECT  11.70 9.54 12.06 9.90 ;
        RECT  20.34 9.54 20.70 9.90 ;
        END
    END rb
    PIN q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  24.60 6.24 26.16 6.72 ;
        RECT  25.32 8.40 25.80 12.36 ;
        RECT  25.56 2.76 26.04 4.56 ;
        RECT  25.68 4.08 26.16 8.88 ;
        END
    END q
    PIN ip
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 7.32 1.32 7.80 ;
        END
    END ip
    PIN ck
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER metal1 ;
        RECT  5.16 6.24 5.64 6.72 ;
        END
    END ck
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.38 0.00 1.86 3.48 ;
        RECT  4.62 0.00 5.10 3.48 ;
        RECT  11.52 0.00 12.00 3.48 ;
        RECT  14.70 0.00 15.18 3.48 ;
        RECT  16.80 0.00 17.28 3.48 ;
        RECT  22.50 0.00 22.98 4.44 ;
        RECT  24.54 0.00 25.02 4.44 ;
        RECT  26.58 0.00 27.06 4.44 ;
        RECT  0.00 0.00 28.08 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.66 10.44 1.14 15.12 ;
        RECT  3.36 10.44 3.84 15.12 ;
        RECT  4.44 10.44 4.92 15.12 ;
        RECT  10.80 10.44 11.28 15.12 ;
        RECT  14.70 10.44 15.18 15.12 ;
        RECT  16.80 10.44 17.28 15.12 ;
        RECT  20.76 10.44 21.24 15.12 ;
        RECT  24.24 9.06 24.72 15.12 ;
        RECT  26.40 9.18 26.88 15.12 ;
        RECT  0.00 13.80 28.08 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  18.60 9.48 19.08 12.24 ;
        RECT  18.12 7.32 18.60 9.96 ;
        RECT  18.12 7.32 25.08 7.80 ;
        RECT  19.20 4.08 19.68 7.80 ;
        RECT  19.20 4.08 20.22 4.56 ;
        RECT  19.74 3.00 20.22 4.56 ;
        RECT  21.54 5.16 24.06 5.64 ;
        RECT  23.58 2.76 24.06 5.64 ;
        RECT  21.54 3.00 22.02 5.64 ;
        RECT  22.44 11.58 23.04 12.18 ;
        RECT  22.50 9.06 22.98 12.18 ;
        RECT  20.22 5.10 20.82 5.70 ;
        RECT  19.68 11.58 20.28 12.18 ;
        RECT  19.74 10.44 20.22 12.18 ;
        RECT  19.14 8.34 19.74 8.94 ;
        RECT  17.76 3.00 19.20 3.48 ;
        RECT  18.06 6.18 18.66 6.78 ;
        RECT  18.12 4.02 18.60 6.78 ;
        RECT  18.06 4.02 18.66 4.62 ;
        RECT  15.72 9.48 16.20 12.12 ;
        RECT  15.96 4.08 16.44 9.96 ;
        RECT  15.90 7.26 16.50 7.86 ;
        RECT  15.90 7.32 17.52 7.80 ;
        RECT  15.72 3.00 16.20 4.56 ;
        RECT  7.92 7.32 8.40 12.24 ;
        RECT  7.92 8.40 14.46 8.88 ;
        RECT  13.98 7.32 14.46 8.88 ;
        RECT  13.98 7.32 15.36 7.80 ;
        RECT  7.80 3.00 8.28 7.80 ;
        RECT  13.50 2.94 14.10 3.54 ;
        RECT  10.56 4.08 12.96 4.56 ;
        RECT  12.48 3.00 12.96 4.56 ;
        RECT  10.56 3.00 11.04 4.56 ;
        RECT  11.76 11.58 12.36 12.18 ;
        RECT  11.82 10.44 12.30 12.18 ;
        RECT  10.50 7.26 11.10 7.86 ;
        RECT  9.42 4.02 10.02 4.62 ;
        RECT  8.88 11.58 9.48 12.18 ;
        RECT  8.94 10.44 9.42 12.18 ;
        RECT  8.76 2.94 9.36 3.54 ;
        RECT  6.84 11.58 7.44 12.18 ;
        RECT  6.90 10.44 7.38 12.18 ;
        RECT  6.72 2.94 7.32 3.54 ;
        RECT  5.52 9.48 6.00 12.12 ;
        RECT  5.52 9.48 6.72 9.96 ;
        RECT  6.24 4.08 6.72 9.96 ;
        RECT  6.18 6.18 6.78 6.78 ;
        RECT  5.64 4.08 6.72 4.56 ;
        RECT  5.64 3.00 6.12 4.56 ;
        RECT  5.10 8.34 5.70 8.94 ;
        RECT  4.02 4.02 4.62 4.62 ;
        RECT  3.36 2.94 3.96 3.54 ;
        RECT  2.34 11.58 2.94 12.18 ;
        RECT  2.40 10.44 2.88 12.18 ;
        RECT  0.42 4.08 2.82 4.56 ;
        RECT  2.34 3.00 2.82 4.56 ;
        RECT  0.42 3.00 0.90 4.56 ;
        LAYER via ;
        RECT  22.56 11.70 22.92 12.06 ;
        RECT  20.34 5.22 20.70 5.58 ;
        RECT  19.80 11.70 20.16 12.06 ;
        RECT  19.26 8.46 19.62 8.82 ;
        RECT  18.18 4.14 18.54 4.50 ;
        RECT  18.18 6.30 18.54 6.66 ;
        RECT  16.02 7.38 16.38 7.74 ;
        RECT  13.62 3.06 13.98 3.42 ;
        RECT  11.88 11.70 12.24 12.06 ;
        RECT  10.62 7.38 10.98 7.74 ;
        RECT  9.54 4.14 9.90 4.50 ;
        RECT  9.00 11.70 9.36 12.06 ;
        RECT  8.88 3.06 9.24 3.42 ;
        RECT  6.96 11.70 7.32 12.06 ;
        RECT  6.84 3.06 7.20 3.42 ;
        RECT  6.30 6.30 6.66 6.66 ;
        RECT  5.22 8.46 5.58 8.82 ;
        RECT  4.14 4.14 4.50 4.50 ;
        RECT  3.48 3.06 3.84 3.42 ;
        RECT  2.46 11.70 2.82 12.06 ;
        LAYER metal2 ;
        RECT  22.44 11.58 23.04 12.18 ;
        RECT  19.68 11.58 20.28 12.18 ;
        RECT  19.68 11.64 23.04 12.12 ;
        RECT  20.22 5.10 20.82 5.70 ;
        RECT  20.28 4.08 20.76 5.70 ;
        RECT  18.06 4.02 18.66 4.62 ;
        RECT  18.06 4.08 20.76 4.56 ;
        RECT  19.14 8.34 19.74 8.94 ;
        RECT  5.10 8.34 5.70 8.94 ;
        RECT  5.10 8.40 19.74 8.88 ;
        RECT  18.06 6.18 18.66 6.78 ;
        RECT  6.18 6.18 6.78 6.78 ;
        RECT  6.18 6.24 18.66 6.72 ;
        RECT  15.90 7.26 16.50 7.86 ;
        RECT  10.50 7.26 11.10 7.86 ;
        RECT  10.50 7.32 16.50 7.80 ;
        RECT  13.50 2.94 14.10 3.54 ;
        RECT  8.76 2.94 9.36 3.54 ;
        RECT  8.76 3.00 14.10 3.48 ;
        RECT  11.76 11.58 12.36 12.18 ;
        RECT  8.88 11.58 9.48 12.18 ;
        RECT  8.88 11.64 12.36 12.12 ;
        RECT  9.42 4.02 10.02 4.62 ;
        RECT  4.02 4.02 4.62 4.62 ;
        RECT  4.02 4.08 10.02 4.56 ;
        RECT  6.84 11.58 7.44 12.18 ;
        RECT  2.34 11.58 2.94 12.18 ;
        RECT  2.34 11.64 7.44 12.12 ;
        RECT  6.72 2.94 7.32 3.54 ;
        RECT  3.36 2.94 3.96 3.54 ;
        RECT  3.36 3.00 7.32 3.48 ;
    END
END drsp_4

MACRO dtrsp_2
    CLASS CORE ;
    FOREIGN dtrsp_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 43.20 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN sm
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal2 ;
        RECT  1.86 8.34 2.46 8.94 ;
        RECT  1.86 8.40 7.86 8.88 ;
        RECT  7.26 8.34 7.86 8.94 ;
        LAYER metal1 ;
        RECT  1.86 8.34 2.46 8.94 ;
        RECT  7.26 8.34 7.86 8.94 ;
        LAYER via ;
        RECT  1.98 8.46 2.34 8.82 ;
        RECT  7.38 8.46 7.74 8.82 ;
        END
    END sm
    PIN sip
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  4.08 6.24 4.56 6.72 ;
        END
    END sip
    PIN s
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal2 ;
        RECT  12.66 5.10 13.26 5.70 ;
        RECT  22.38 5.10 22.98 5.70 ;
        RECT  12.66 5.16 32.64 5.64 ;
        RECT  32.16 5.16 32.64 6.72 ;
        RECT  36.48 5.10 36.96 6.72 ;
        RECT  32.16 6.24 36.96 6.72 ;
        RECT  36.42 5.10 37.02 5.70 ;
        LAYER metal1 ;
        RECT  12.66 5.10 13.26 5.70 ;
        RECT  22.38 5.10 22.98 5.70 ;
        RECT  36.42 5.10 37.02 5.70 ;
        LAYER via ;
        RECT  12.78 5.22 13.14 5.58 ;
        RECT  22.50 5.22 22.86 5.58 ;
        RECT  36.54 5.22 36.90 5.58 ;
        END
    END s
    PIN rb
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal2 ;
        RECT  13.74 9.42 14.34 10.02 ;
        RECT  24.54 9.42 25.14 10.02 ;
        RECT  13.74 9.48 34.86 9.96 ;
        RECT  34.26 9.42 34.86 10.02 ;
        LAYER metal1 ;
        RECT  13.74 9.42 14.34 10.02 ;
        RECT  24.54 9.42 25.14 10.02 ;
        RECT  34.26 9.42 34.86 10.02 ;
        LAYER via ;
        RECT  13.86 9.54 14.22 9.90 ;
        RECT  24.66 9.54 25.02 9.90 ;
        RECT  34.38 9.54 34.74 9.90 ;
        END
    END rb
    PIN q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  39.72 3.00 40.20 6.72 ;
        RECT  38.64 6.24 41.28 6.72 ;
        RECT  39.72 3.00 40.80 3.48 ;
        RECT  40.32 8.40 40.80 12.30 ;
        RECT  40.80 6.24 41.28 8.88 ;
        END
    END q
    PIN ip
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  6.24 7.32 6.72 7.80 ;
        END
    END ip
    PIN ck
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER metal1 ;
        RECT  15.96 6.24 16.44 6.72 ;
        END
    END ck
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.58 0.00 3.06 3.48 ;
        RECT  7.86 0.00 8.34 3.48 ;
        RECT  12.18 0.00 12.66 3.48 ;
        RECT  15.72 0.00 16.20 3.48 ;
        RECT  23.40 0.00 23.88 3.48 ;
        RECT  26.88 0.00 27.36 3.48 ;
        RECT  29.52 0.00 30.00 3.48 ;
        RECT  36.54 0.00 37.02 3.48 ;
        RECT  38.76 0.00 39.24 3.48 ;
        RECT  41.58 0.00 42.06 3.48 ;
        RECT  0.00 0.00 43.20 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.64 10.62 3.12 15.12 ;
        RECT  7.92 10.62 8.40 15.12 ;
        RECT  11.10 10.62 11.58 15.12 ;
        RECT  14.34 10.62 14.82 15.12 ;
        RECT  15.66 10.62 16.14 15.12 ;
        RECT  22.92 10.62 23.40 15.12 ;
        RECT  26.64 10.62 27.12 15.12 ;
        RECT  29.52 10.62 30.00 15.12 ;
        RECT  33.96 10.62 34.44 15.12 ;
        RECT  38.76 10.62 39.24 15.12 ;
        RECT  41.64 10.62 42.12 15.12 ;
        RECT  0.00 13.80 43.20 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  40.74 5.10 41.34 5.70 ;
        RECT  31.68 7.32 32.16 12.30 ;
        RECT  39.66 7.26 40.26 7.86 ;
        RECT  31.68 7.32 40.26 7.80 ;
        RECT  33.24 3.00 33.72 7.80 ;
        RECT  35.52 4.14 38.10 4.62 ;
        RECT  37.62 3.00 38.10 4.62 ;
        RECT  35.52 3.00 36.00 4.62 ;
        RECT  36.54 10.62 37.02 12.30 ;
        RECT  36.48 11.58 37.08 12.18 ;
        RECT  34.26 5.10 34.86 5.70 ;
        RECT  33.18 8.34 33.78 8.94 ;
        RECT  32.94 10.62 33.42 12.30 ;
        RECT  32.88 11.58 33.48 12.18 ;
        RECT  30.60 3.00 32.46 3.48 ;
        RECT  31.02 6.18 31.62 6.78 ;
        RECT  31.08 4.02 31.56 6.78 ;
        RECT  31.02 4.02 31.62 4.62 ;
        RECT  28.26 3.00 28.74 12.30 ;
        RECT  28.26 7.26 29.46 7.86 ;
        RECT  28.26 7.32 30.48 7.80 ;
        RECT  19.44 3.00 19.92 12.30 ;
        RECT  19.44 8.40 25.08 8.88 ;
        RECT  24.60 7.32 25.08 8.88 ;
        RECT  24.60 7.32 27.24 7.80 ;
        RECT  25.62 2.94 26.22 3.54 ;
        RECT  22.38 4.02 24.96 4.50 ;
        RECT  24.48 2.82 24.96 4.50 ;
        RECT  22.38 2.82 22.86 4.50 ;
        RECT  24.30 10.62 24.78 12.30 ;
        RECT  24.24 11.58 24.84 12.18 ;
        RECT  22.38 7.26 22.98 7.86 ;
        RECT  21.30 4.02 21.90 4.62 ;
        RECT  20.88 2.94 21.48 3.54 ;
        RECT  20.70 10.62 21.18 12.30 ;
        RECT  20.64 11.58 21.24 12.18 ;
        RECT  18.30 2.94 18.90 3.54 ;
        RECT  18.30 10.62 18.78 12.30 ;
        RECT  18.24 11.58 18.84 12.18 ;
        RECT  17.04 3.00 17.52 12.30 ;
        RECT  16.98 6.18 17.58 6.78 ;
        RECT  15.90 4.02 16.50 4.62 ;
        RECT  15.90 8.34 16.50 8.94 ;
        RECT  14.46 2.94 15.06 3.54 ;
        RECT  13.20 10.62 13.68 12.30 ;
        RECT  13.14 11.58 13.74 12.18 ;
        RECT  11.10 4.02 13.68 4.50 ;
        RECT  13.20 3.00 13.68 4.50 ;
        RECT  11.10 3.00 11.58 4.50 ;
        RECT  9.60 8.40 10.08 12.30 ;
        RECT  9.60 8.40 11.04 8.88 ;
        RECT  10.56 5.16 11.04 8.88 ;
        RECT  10.56 6.24 12.12 6.72 ;
        RECT  9.60 5.16 11.04 5.64 ;
        RECT  9.60 3.00 10.08 5.64 ;
        RECT  5.34 3.00 5.82 12.30 ;
        RECT  5.34 6.24 9.42 6.72 ;
        RECT  7.26 5.10 7.86 5.70 ;
        RECT  0.90 3.00 1.38 12.30 ;
        RECT  2.94 5.10 3.54 5.70 ;
        RECT  0.90 5.16 3.54 5.64 ;
        LAYER via ;
        RECT  40.86 5.22 41.22 5.58 ;
        RECT  39.78 7.38 40.14 7.74 ;
        RECT  36.60 11.70 36.96 12.06 ;
        RECT  34.38 5.22 34.74 5.58 ;
        RECT  33.30 8.46 33.66 8.82 ;
        RECT  33.00 11.70 33.36 12.06 ;
        RECT  31.14 4.14 31.50 4.50 ;
        RECT  31.14 6.30 31.50 6.66 ;
        RECT  28.98 7.38 29.34 7.74 ;
        RECT  25.74 3.06 26.10 3.42 ;
        RECT  24.36 11.70 24.72 12.06 ;
        RECT  22.50 7.38 22.86 7.74 ;
        RECT  21.42 4.14 21.78 4.50 ;
        RECT  21.00 3.06 21.36 3.42 ;
        RECT  20.76 11.70 21.12 12.06 ;
        RECT  18.42 3.06 18.78 3.42 ;
        RECT  18.36 11.70 18.72 12.06 ;
        RECT  17.10 6.30 17.46 6.66 ;
        RECT  16.02 4.14 16.38 4.50 ;
        RECT  16.02 8.46 16.38 8.82 ;
        RECT  14.58 3.06 14.94 3.42 ;
        RECT  13.26 11.70 13.62 12.06 ;
        RECT  7.38 5.22 7.74 5.58 ;
        RECT  3.06 5.22 3.42 5.58 ;
        LAYER metal2 ;
        RECT  39.66 7.26 40.26 7.86 ;
        RECT  39.72 5.16 40.20 7.86 ;
        RECT  40.74 5.10 41.34 5.70 ;
        RECT  39.72 5.16 41.34 5.64 ;
        RECT  36.48 11.58 37.08 12.18 ;
        RECT  32.88 11.58 33.48 12.18 ;
        RECT  32.88 11.64 37.08 12.12 ;
        RECT  34.26 5.10 34.86 5.70 ;
        RECT  34.32 4.08 34.80 5.70 ;
        RECT  31.02 4.02 31.62 4.62 ;
        RECT  31.02 4.08 34.80 4.56 ;
        RECT  33.18 8.34 33.78 8.94 ;
        RECT  15.90 8.34 16.50 8.94 ;
        RECT  15.90 8.40 33.78 8.88 ;
        RECT  31.02 6.18 31.62 6.78 ;
        RECT  16.98 6.18 17.58 6.78 ;
        RECT  16.98 6.24 31.62 6.72 ;
        RECT  28.86 7.26 29.46 7.86 ;
        RECT  22.38 7.26 22.98 7.86 ;
        RECT  22.38 7.32 29.46 7.80 ;
        RECT  25.62 2.94 26.22 3.54 ;
        RECT  20.88 2.94 21.48 3.54 ;
        RECT  20.88 3.00 26.22 3.48 ;
        RECT  24.24 11.58 24.84 12.18 ;
        RECT  20.64 11.58 21.24 12.18 ;
        RECT  20.64 11.64 24.84 12.12 ;
        RECT  21.30 4.02 21.90 4.62 ;
        RECT  15.90 4.02 16.50 4.62 ;
        RECT  15.90 4.08 21.90 4.56 ;
        RECT  18.30 2.94 18.90 3.54 ;
        RECT  14.46 2.94 15.06 3.54 ;
        RECT  14.46 3.00 18.90 3.48 ;
        RECT  18.24 11.58 18.84 12.18 ;
        RECT  13.14 11.58 13.74 12.18 ;
        RECT  13.14 11.64 18.84 12.12 ;
        RECT  7.26 5.10 7.86 5.70 ;
        RECT  2.94 5.10 3.54 5.70 ;
        RECT  2.94 5.16 7.86 5.64 ;
    END
END dtrsp_2

MACRO filler
    CLASS CORE ;
    FOREIGN filler 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 1.08 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.00 0.00 1.08 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.00 13.80 1.08 15.12 ;
        END
    END vdd
END filler

MACRO fulladder
    CLASS CORE ;
    FOREIGN fulladder 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.76 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN s
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  22.44 2.94 22.92 12.36 ;
        END
    END s
    PIN co
        DIRECTION OUTPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  10.02 3.00 10.50 4.56 ;
        RECT  10.02 9.48 10.50 12.36 ;
        RECT  10.02 4.08 11.04 4.56 ;
        RECT  10.56 4.08 11.04 9.96 ;
        RECT  10.02 9.48 11.04 9.96 ;
        END
    END co
    PIN ci
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal2 ;
        RECT  5.10 6.18 5.70 6.78 ;
        RECT  13.74 6.18 14.34 6.78 ;
        RECT  5.10 6.24 20.82 6.72 ;
        RECT  20.22 6.18 20.82 6.78 ;
        LAYER metal1 ;
        RECT  5.10 6.18 5.70 6.78 ;
        RECT  13.74 6.18 14.34 6.78 ;
        RECT  20.22 6.18 20.82 6.78 ;
        LAYER via ;
        RECT  5.22 6.30 5.58 6.66 ;
        RECT  13.86 6.30 14.22 6.66 ;
        RECT  20.34 6.30 20.70 6.66 ;
        END
    END ci
    PIN b
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal2 ;
        RECT  2.94 7.26 3.54 7.86 ;
        RECT  8.34 7.26 8.94 7.86 ;
        RECT  12.66 7.26 13.26 7.86 ;
        RECT  2.94 7.32 18.66 7.80 ;
        RECT  18.06 7.26 18.66 7.86 ;
        LAYER metal1 ;
        RECT  2.94 7.26 3.54 7.86 ;
        RECT  8.34 7.26 8.94 7.86 ;
        RECT  12.66 7.26 13.26 7.86 ;
        RECT  18.06 7.26 18.66 7.86 ;
        LAYER via ;
        RECT  3.06 7.38 3.42 7.74 ;
        RECT  8.46 7.38 8.82 7.74 ;
        RECT  12.78 7.38 13.14 7.74 ;
        RECT  18.18 7.38 18.54 7.74 ;
        END
    END b
    PIN a
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal2 ;
        RECT  0.78 8.34 1.38 8.94 ;
        RECT  6.18 8.34 6.78 8.94 ;
        RECT  11.58 8.34 12.18 8.94 ;
        RECT  0.78 8.40 17.58 8.88 ;
        RECT  16.98 8.34 17.58 8.94 ;
        LAYER metal1 ;
        RECT  0.78 8.34 1.38 8.94 ;
        RECT  6.18 8.34 6.78 8.94 ;
        RECT  11.58 8.34 12.18 8.94 ;
        RECT  16.98 8.34 17.58 8.94 ;
        LAYER via ;
        RECT  0.90 8.46 1.26 8.82 ;
        RECT  6.30 8.46 6.66 8.82 ;
        RECT  11.70 8.46 12.06 8.82 ;
        RECT  17.10 8.46 17.46 8.82 ;
        END
    END a
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.90 0.00 1.38 3.48 ;
        RECT  5.94 0.00 6.42 3.48 ;
        RECT  7.98 0.00 8.46 3.48 ;
        RECT  9.00 0.00 9.48 3.48 ;
        RECT  10.98 0.00 11.46 3.48 ;
        RECT  18.12 0.00 18.60 3.48 ;
        RECT  20.16 0.00 20.64 3.48 ;
        RECT  21.42 0.00 21.90 3.48 ;
        RECT  0.00 0.00 23.76 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.90 10.68 1.38 15.12 ;
        RECT  2.94 10.68 3.42 15.12 ;
        RECT  9.00 10.68 9.48 15.12 ;
        RECT  10.98 10.68 11.46 15.12 ;
        RECT  13.02 10.68 13.50 15.12 ;
        RECT  21.42 10.68 21.90 15.12 ;
        RECT  0.00 13.80 23.76 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  20.16 9.48 20.64 12.36 ;
        RECT  15.12 3.00 15.60 12.36 ;
        RECT  20.16 9.48 21.84 9.96 ;
        RECT  21.36 5.16 21.84 9.96 ;
        RECT  15.12 5.16 21.84 5.64 ;
        RECT  14.04 3.00 15.60 3.48 ;
        RECT  19.08 2.94 19.68 3.54 ;
        RECT  17.10 2.94 17.70 3.54 ;
        RECT  16.14 3.00 17.70 3.48 ;
        RECT  16.98 9.42 17.58 10.02 ;
        RECT  17.10 10.68 17.58 12.36 ;
        RECT  16.14 10.68 16.62 12.36 ;
        RECT  16.08 11.58 16.68 12.18 ;
        RECT  16.08 11.64 17.58 12.12 ;
        RECT  14.04 10.68 14.52 12.36 ;
        RECT  13.98 11.58 14.58 12.18 ;
        RECT  12.00 10.68 12.48 12.36 ;
        RECT  11.94 11.58 12.54 12.18 ;
        RECT  7.98 9.48 8.46 12.36 ;
        RECT  3.90 3.00 4.38 12.36 ;
        RECT  8.34 9.42 8.94 10.02 ;
        RECT  3.90 9.48 9.18 9.96 ;
        RECT  2.94 3.00 4.38 3.48 ;
        RECT  6.90 2.94 7.50 3.54 ;
        RECT  5.94 10.62 6.42 12.30 ;
        RECT  4.92 10.62 5.40 12.30 ;
        RECT  4.86 11.58 5.46 12.18 ;
        RECT  4.86 11.64 6.42 12.12 ;
        RECT  4.86 2.94 5.46 3.54 ;
        RECT  1.92 10.62 2.40 12.30 ;
        RECT  1.86 11.58 2.46 12.18 ;
        LAYER via ;
        RECT  19.20 3.06 19.56 3.42 ;
        RECT  17.22 3.06 17.58 3.42 ;
        RECT  17.10 9.54 17.46 9.90 ;
        RECT  16.20 11.70 16.56 12.06 ;
        RECT  14.10 11.70 14.46 12.06 ;
        RECT  12.06 11.70 12.42 12.06 ;
        RECT  8.46 9.54 8.82 9.90 ;
        RECT  7.02 3.06 7.38 3.42 ;
        RECT  4.98 3.06 5.34 3.42 ;
        RECT  4.98 11.70 5.34 12.06 ;
        RECT  1.98 11.70 2.34 12.06 ;
        LAYER metal2 ;
        RECT  19.08 2.94 19.68 3.54 ;
        RECT  17.10 2.94 17.70 3.54 ;
        RECT  17.10 3.00 19.68 3.48 ;
        RECT  16.98 9.42 17.58 10.02 ;
        RECT  8.34 9.42 8.94 10.02 ;
        RECT  8.28 9.48 17.58 9.96 ;
        RECT  16.08 11.58 16.68 12.18 ;
        RECT  13.98 11.58 14.58 12.18 ;
        RECT  11.94 11.58 12.54 12.18 ;
        RECT  11.94 11.64 16.68 12.12 ;
        RECT  6.90 2.94 7.50 3.54 ;
        RECT  4.86 2.94 5.46 3.54 ;
        RECT  4.86 3.00 7.50 3.48 ;
        RECT  4.86 11.58 5.46 12.18 ;
        RECT  1.86 11.58 2.46 12.18 ;
        RECT  1.86 11.64 5.46 12.12 ;
    END
END fulladder

MACRO inv_1
    CLASS CORE ;
    FOREIGN inv_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 3.24 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.92 3.00 2.40 12.36 ;
        END
    END op
    PIN ip
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 7.32 1.32 7.80 ;
        END
    END ip
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.90 0.00 1.38 3.48 ;
        RECT  0.00 0.00 3.24 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.90 10.68 1.38 15.12 ;
        RECT  0.00 13.80 3.24 15.12 ;
        END
    END vdd
END inv_1

MACRO inv_2
    CLASS CORE ;
    FOREIGN inv_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 3.24 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.92 2.76 2.40 12.36 ;
        END
    END op
    PIN ip
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 6.24 1.32 6.72 ;
        END
    END ip
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.90 0.00 1.38 4.44 ;
        RECT  0.00 0.00 3.24 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.90 9.00 1.38 15.12 ;
        RECT  0.00 13.80 3.24 15.12 ;
        END
    END vdd
END inv_2

MACRO inv_4
    CLASS CORE ;
    FOREIGN inv_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 3.24 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.76 1.92 5.64 ;
        RECT  1.44 7.32 1.92 12.36 ;
        RECT  1.92 5.16 2.40 7.80 ;
        END
    END op
    PIN ip
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 6.24 1.32 6.72 ;
        END
    END ip
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.42 0.00 0.90 4.44 ;
        RECT  2.46 0.00 2.94 4.44 ;
        RECT  0.00 0.00 3.24 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.42 9.00 0.90 15.12 ;
        RECT  2.40 9.00 2.88 15.12 ;
        RECT  0.00 13.80 3.24 15.12 ;
        END
    END vdd
END inv_4

MACRO invzp_1
    CLASS CORE ;
    FOREIGN invzp_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.40 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.72 3.00 4.20 4.56 ;
        RECT  3.72 10.56 4.20 12.36 ;
        RECT  4.08 4.08 4.56 11.04 ;
        END
    END op
    PIN ip
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  1.92 6.24 2.40 6.72 ;
        END
    END ip
    PIN c
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  1.92 7.32 3.48 7.80 ;
        RECT  3.00 7.32 3.48 9.96 ;
        END
    END c
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.92 0.00 2.40 3.48 ;
        RECT  0.00 0.00 5.40 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.92 10.92 2.40 15.12 ;
        RECT  0.00 13.80 5.40 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  0.60 3.00 1.08 12.36 ;
        RECT  0.60 5.16 3.48 5.64 ;
    END
END invzp_1

MACRO invzp_2
    CLASS CORE ;
    FOREIGN invzp_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.48 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.26 2.76 4.74 4.44 ;
        RECT  4.26 8.40 4.74 12.36 ;
        RECT  4.26 3.96 5.64 4.44 ;
        RECT  5.16 3.96 5.64 8.88 ;
        RECT  4.26 8.40 5.64 8.88 ;
        END
    END op
    PIN ip
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  3.00 6.24 3.48 6.72 ;
        END
    END ip
    PIN c
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  1.92 7.32 4.56 7.80 ;
        END
    END c
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.46 0.00 2.94 4.44 ;
        RECT  0.00 0.00 6.48 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.46 9.00 2.94 15.12 ;
        RECT  0.00 13.80 6.48 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  1.14 8.40 1.62 12.36 ;
        RECT  0.84 4.08 1.32 8.88 ;
        RECT  0.84 5.16 4.56 5.64 ;
        RECT  1.14 2.76 1.62 4.56 ;
    END
END invzp_2

MACRO invzp_4
    CLASS CORE ;
    FOREIGN invzp_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.48 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.78 2.76 4.26 4.68 ;
        RECT  3.90 8.40 4.38 12.36 ;
        RECT  3.78 4.20 5.64 4.68 ;
        RECT  5.16 4.20 5.64 8.88 ;
        RECT  3.90 8.40 5.64 8.88 ;
        END
    END op
    PIN ip
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  4.08 6.24 4.56 6.72 ;
        END
    END ip
    PIN c
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  1.92 6.24 2.40 7.80 ;
        RECT  1.92 7.32 4.56 7.80 ;
        END
    END c
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.98 0.00 2.46 4.32 ;
        RECT  5.58 0.00 6.06 3.84 ;
        RECT  0.00 0.00 6.48 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.10 9.00 2.58 15.12 ;
        RECT  5.70 9.24 6.18 15.12 ;
        RECT  0.00 13.80 6.48 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  0.78 8.40 1.26 12.36 ;
        RECT  0.48 4.08 0.96 8.88 ;
        RECT  0.48 5.16 4.56 5.64 ;
        RECT  0.78 2.82 1.26 4.56 ;
    END
END invzp_4

MACRO jkrp_2
    CLASS CORE ;
    FOREIGN jkrp_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 35.64 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN rb
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal2 ;
        RECT  21.30 7.26 21.90 7.86 ;
        RECT  21.30 7.32 27.30 7.80 ;
        RECT  26.70 7.26 27.30 7.86 ;
        LAYER metal1 ;
        RECT  21.30 7.26 21.90 7.86 ;
        RECT  26.70 7.26 27.30 7.86 ;
        LAYER via ;
        RECT  21.42 7.38 21.78 7.74 ;
        RECT  26.82 7.38 27.18 7.74 ;
        END
    END rb
    PIN qb
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  32.88 2.76 33.36 12.36 ;
        RECT  32.88 6.24 33.72 7.80 ;
        END
    END qb
    PIN q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  34.32 7.32 35.34 7.80 ;
        RECT  34.86 2.76 35.34 12.36 ;
        END
    END q
    PIN k
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  5.16 8.40 5.64 8.88 ;
        END
    END k
    PIN j
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 7.32 1.32 7.80 ;
        END
    END j
    PIN ck
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER metal1 ;
        RECT  10.14 6.30 10.62 6.78 ;
        END
    END ck
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.66 0.00 1.14 3.66 ;
        RECT  2.76 0.00 3.24 3.66 ;
        RECT  6.84 0.00 7.32 3.66 ;
        RECT  10.14 0.00 10.62 3.66 ;
        RECT  12.12 0.00 12.60 3.66 ;
        RECT  16.80 0.00 17.28 3.66 ;
        RECT  19.14 0.00 19.62 3.66 ;
        RECT  26.88 0.00 27.36 3.66 ;
        RECT  29.88 0.00 30.36 3.66 ;
        RECT  31.86 0.00 32.34 4.44 ;
        RECT  33.84 0.00 34.32 4.44 ;
        RECT  0.00 0.00 35.64 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.66 10.68 1.14 15.12 ;
        RECT  3.78 10.68 4.26 15.12 ;
        RECT  10.14 10.68 10.62 15.12 ;
        RECT  12.12 10.68 12.60 15.12 ;
        RECT  16.80 10.68 17.28 15.12 ;
        RECT  19.14 10.68 19.62 15.12 ;
        RECT  21.18 10.68 21.66 15.12 ;
        RECT  26.88 10.68 27.36 15.12 ;
        RECT  28.92 10.68 29.40 15.12 ;
        RECT  29.88 10.68 30.36 15.12 ;
        RECT  31.86 9.00 32.34 15.12 ;
        RECT  33.84 9.00 34.32 15.12 ;
        RECT  0.00 13.80 35.64 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  33.78 5.10 34.38 5.70 ;
        RECT  30.90 2.82 31.38 12.36 ;
        RECT  29.22 9.54 31.38 10.02 ;
        RECT  30.84 7.44 32.34 7.92 ;
        RECT  30.84 4.02 31.44 4.62 ;
        RECT  29.58 6.18 30.18 6.78 ;
        RECT  27.90 5.10 28.38 12.36 ;
        RECT  25.56 2.82 26.04 12.36 ;
        RECT  25.56 8.40 28.38 8.88 ;
        RECT  27.84 5.10 28.44 5.70 ;
        RECT  27.84 5.16 29.40 5.64 ;
        RECT  28.92 2.82 29.40 5.64 ;
        RECT  26.58 9.42 27.30 10.02 ;
        RECT  24.54 2.82 25.02 12.36 ;
        RECT  23.52 2.82 24.00 12.36 ;
        RECT  23.52 7.32 25.02 7.80 ;
        RECT  23.46 6.18 24.06 6.78 ;
        RECT  22.50 2.82 22.98 12.36 ;
        RECT  20.16 5.28 20.64 12.36 ;
        RECT  18.78 8.40 20.64 8.88 ;
        RECT  20.16 5.28 21.66 5.76 ;
        RECT  21.18 2.82 21.66 5.76 ;
        RECT  21.18 5.10 22.98 5.58 ;
        RECT  21.30 6.18 22.02 6.78 ;
        RECT  21.30 8.34 22.02 8.94 ;
        RECT  19.02 7.26 19.62 7.86 ;
        RECT  17.82 2.82 18.30 12.36 ;
        RECT  15.48 2.82 15.96 12.36 ;
        RECT  15.48 9.48 18.30 9.96 ;
        RECT  16.44 8.34 17.04 8.94 ;
        RECT  14.46 2.82 14.94 12.36 ;
        RECT  14.40 7.26 15.00 7.86 ;
        RECT  13.14 5.76 13.62 12.36 ;
        RECT  13.08 9.42 13.68 10.02 ;
        RECT  13.08 6.18 13.68 6.78 ;
        RECT  13.50 4.20 13.98 6.24 ;
        RECT  13.14 2.82 13.62 4.68 ;
        RECT  11.16 2.82 11.64 12.36 ;
        RECT  11.16 8.34 12.18 8.94 ;
        RECT  11.16 7.32 12.60 7.80 ;
        RECT  9.78 4.68 11.64 5.16 ;
        RECT  9.78 9.42 10.50 10.02 ;
        RECT  8.94 2.82 9.42 12.36 ;
        RECT  8.88 7.26 9.48 7.86 ;
        RECT  7.92 2.82 8.40 12.36 ;
        RECT  5.88 9.54 6.36 12.36 ;
        RECT  5.88 9.54 8.40 10.02 ;
        RECT  4.80 6.30 8.40 6.78 ;
        RECT  4.80 2.82 5.28 6.78 ;
        RECT  6.78 4.02 7.38 4.62 ;
        RECT  6.84 10.68 7.32 12.36 ;
        RECT  6.78 11.58 7.38 12.18 ;
        RECT  4.80 10.68 5.28 12.36 ;
        RECT  4.74 11.58 5.34 12.18 ;
        RECT  1.68 8.40 2.16 12.36 ;
        RECT  1.92 4.08 2.40 10.02 ;
        RECT  1.92 7.32 4.80 7.80 ;
        RECT  1.68 3.00 2.16 5.64 ;
        RECT  2.94 5.10 3.54 5.70 ;
        RECT  2.76 10.68 3.24 12.36 ;
        RECT  2.70 11.58 3.30 12.18 ;
        LAYER via ;
        RECT  33.90 5.22 34.26 5.58 ;
        RECT  30.96 4.14 31.32 4.50 ;
        RECT  29.70 6.30 30.06 6.66 ;
        RECT  27.96 5.22 28.32 5.58 ;
        RECT  26.82 9.54 27.18 9.90 ;
        RECT  23.58 6.30 23.94 6.66 ;
        RECT  21.42 6.30 21.78 6.66 ;
        RECT  21.42 8.46 21.78 8.82 ;
        RECT  19.14 7.38 19.50 7.74 ;
        RECT  16.56 8.46 16.92 8.82 ;
        RECT  14.52 7.38 14.88 7.74 ;
        RECT  13.20 6.30 13.56 6.66 ;
        RECT  13.20 9.54 13.56 9.90 ;
        RECT  11.70 8.46 12.06 8.82 ;
        RECT  10.02 9.54 10.38 9.90 ;
        RECT  9.00 7.38 9.36 7.74 ;
        RECT  6.90 4.14 7.26 4.50 ;
        RECT  6.90 11.70 7.26 12.06 ;
        RECT  4.86 11.70 5.22 12.06 ;
        RECT  3.06 5.22 3.42 5.58 ;
        RECT  2.82 11.70 3.18 12.06 ;
        LAYER metal2 ;
        RECT  33.78 5.10 34.38 5.70 ;
        RECT  27.84 5.10 28.44 5.70 ;
        RECT  2.94 5.10 3.54 5.70 ;
        RECT  2.94 5.16 34.38 5.64 ;
        RECT  30.84 4.02 31.44 4.62 ;
        RECT  6.78 4.02 7.38 4.62 ;
        RECT  6.78 4.08 31.44 4.56 ;
        RECT  29.58 6.18 30.18 6.78 ;
        RECT  23.46 6.18 24.06 6.78 ;
        RECT  23.46 6.24 30.18 6.72 ;
        RECT  26.58 9.42 27.30 10.02 ;
        RECT  13.08 9.42 13.68 10.02 ;
        RECT  9.90 9.42 10.50 10.02 ;
        RECT  9.90 9.48 27.30 9.96 ;
        RECT  21.30 6.18 21.90 6.78 ;
        RECT  13.08 6.18 13.68 6.78 ;
        RECT  13.08 6.24 21.90 6.72 ;
        RECT  21.30 8.34 21.90 8.94 ;
        RECT  16.44 8.34 17.04 8.94 ;
        RECT  11.58 8.34 12.18 8.94 ;
        RECT  11.58 8.40 21.90 8.88 ;
        RECT  19.02 7.26 19.62 7.86 ;
        RECT  14.40 7.26 15.00 7.86 ;
        RECT  8.88 7.26 9.48 7.86 ;
        RECT  8.88 7.32 19.62 7.80 ;
        RECT  6.78 11.58 7.38 12.18 ;
        RECT  4.74 11.58 5.34 12.18 ;
        RECT  2.70 11.58 3.30 12.18 ;
        RECT  2.70 11.64 7.38 12.12 ;
    END
END jkrp_2

MACRO lp_1
    CLASS CORE ;
    FOREIGN lp_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.72 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.56 3.00 8.04 5.64 ;
        RECT  7.56 9.48 8.04 12.36 ;
        RECT  6.24 5.16 8.88 5.64 ;
        RECT  8.40 5.16 8.88 9.96 ;
        RECT  7.56 9.48 8.88 9.96 ;
        END
    END q
    PIN ip
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  3.00 6.24 3.48 6.72 ;
        END
    END ip
    PIN ck
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER metal1 ;
        RECT  1.92 5.16 4.56 5.64 ;
        END
    END ck
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.70 0.00 3.18 3.48 ;
        RECT  6.48 0.00 6.96 3.48 ;
        RECT  8.70 0.00 9.18 3.48 ;
        RECT  0.00 0.00 9.72 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.70 10.68 3.18 15.12 ;
        RECT  6.54 10.68 7.02 15.12 ;
        RECT  8.64 10.68 9.12 15.12 ;
        RECT  0.00 13.80 9.72 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  4.62 10.32 5.10 12.36 ;
        RECT  4.62 10.32 6.12 10.80 ;
        RECT  5.64 8.40 6.12 10.80 ;
        RECT  5.64 8.40 6.72 8.88 ;
        RECT  6.24 6.24 6.72 8.88 ;
        RECT  5.16 6.24 7.80 6.72 ;
        RECT  5.16 4.08 5.64 6.72 ;
        RECT  4.50 4.08 5.64 4.56 ;
        RECT  4.50 3.00 4.98 4.56 ;
        RECT  1.92 7.32 5.64 7.80 ;
        RECT  1.62 9.48 2.10 12.36 ;
        RECT  0.84 9.48 4.56 9.96 ;
        RECT  0.84 4.08 1.32 9.96 ;
        RECT  0.84 4.08 2.10 4.56 ;
        RECT  1.62 3.00 2.10 4.56 ;
    END
END lp_1

MACRO lp_2
    CLASS CORE ;
    FOREIGN lp_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.72 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.56 2.76 8.04 5.64 ;
        RECT  7.56 8.40 8.04 12.36 ;
        RECT  6.24 5.16 8.88 5.64 ;
        RECT  8.40 5.16 8.88 8.88 ;
        RECT  7.56 8.40 8.88 8.88 ;
        END
    END q
    PIN ip
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  3.00 6.24 3.48 6.72 ;
        END
    END ip
    PIN ck
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER metal1 ;
        RECT  1.92 5.16 4.56 5.64 ;
        END
    END ck
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.70 0.00 3.18 4.32 ;
        RECT  6.48 0.00 6.96 4.32 ;
        RECT  8.70 0.00 9.18 4.32 ;
        RECT  0.00 0.00 9.72 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.70 9.24 3.18 15.12 ;
        RECT  6.54 9.24 7.02 15.12 ;
        RECT  8.64 9.24 9.12 15.12 ;
        RECT  0.00 13.80 9.72 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  4.62 9.24 5.10 12.36 ;
        RECT  4.62 9.24 6.12 9.72 ;
        RECT  5.64 8.40 6.12 9.72 ;
        RECT  5.64 8.40 6.96 8.88 ;
        RECT  6.48 6.24 6.96 8.88 ;
        RECT  5.16 6.24 7.80 6.72 ;
        RECT  5.16 4.08 5.64 6.72 ;
        RECT  4.50 4.08 5.64 4.56 ;
        RECT  4.50 2.76 4.98 4.56 ;
        RECT  1.92 7.32 5.64 7.80 ;
        RECT  1.62 8.40 2.10 12.36 ;
        RECT  0.84 8.40 4.56 8.88 ;
        RECT  0.84 4.08 1.32 8.88 ;
        RECT  0.84 4.08 2.10 4.56 ;
        RECT  1.62 2.76 2.10 4.56 ;
    END
END lp_2

MACRO lrp_1
    CLASS CORE ;
    FOREIGN lrp_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.04 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN rb
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal2 ;
        RECT  1.86 8.34 2.46 8.94 ;
        RECT  1.86 8.40 10.02 8.88 ;
        RECT  9.42 8.34 10.02 8.94 ;
        LAYER metal1 ;
        RECT  1.86 8.34 2.46 8.94 ;
        RECT  9.42 8.34 10.02 8.94 ;
        LAYER via ;
        RECT  1.98 8.46 2.34 8.82 ;
        RECT  9.54 8.46 9.90 8.82 ;
        END
    END rb
    PIN q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.40 6.24 13.20 6.72 ;
        RECT  12.72 4.08 13.20 9.96 ;
        RECT  12.96 3.00 13.44 4.56 ;
        RECT  12.96 9.48 13.44 12.12 ;
        END
    END q
    PIN ip
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 6.24 1.32 6.72 ;
        END
    END ip
    PIN ck
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER metal2 ;
        RECT  4.02 6.18 4.62 6.78 ;
        RECT  4.02 6.24 7.86 6.72 ;
        RECT  7.26 6.18 7.86 6.78 ;
        LAYER metal1 ;
        RECT  4.08 6.18 4.56 7.80 ;
        RECT  4.02 6.18 4.62 6.78 ;
        RECT  7.26 6.18 7.86 6.78 ;
        LAYER via ;
        RECT  4.14 6.30 4.50 6.66 ;
        RECT  7.38 6.30 7.74 6.66 ;
        END
    END ck
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.60 0.00 1.08 3.48 ;
        RECT  3.54 0.00 4.02 3.48 ;
        RECT  8.94 0.00 9.42 3.48 ;
        RECT  11.94 0.00 12.42 3.48 ;
        RECT  0.00 0.00 14.04 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.30 10.44 0.78 15.12 ;
        RECT  2.28 10.44 2.76 15.12 ;
        RECT  3.36 10.44 3.84 15.12 ;
        RECT  8.88 10.44 9.36 15.12 ;
        RECT  11.94 10.44 12.42 15.12 ;
        RECT  0.00 13.80 14.04 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  6.84 9.48 7.32 12.12 ;
        RECT  6.24 9.48 7.32 9.96 ;
        RECT  6.24 5.16 6.72 9.96 ;
        RECT  6.24 7.32 12.12 7.80 ;
        RECT  6.72 3.00 7.20 5.64 ;
        RECT  7.74 4.08 11.34 4.56 ;
        RECT  10.86 3.00 11.34 4.56 ;
        RECT  7.74 3.00 8.22 4.56 ;
        RECT  9.96 9.48 10.44 12.12 ;
        RECT  7.86 9.48 8.34 12.12 ;
        RECT  7.86 9.48 10.44 9.96 ;
        RECT  5.76 11.58 6.36 12.18 ;
        RECT  5.82 10.44 6.30 12.18 ;
        RECT  5.64 2.94 6.24 3.54 ;
        RECT  4.44 9.48 4.92 12.12 ;
        RECT  4.44 9.48 5.64 9.96 ;
        RECT  5.16 4.08 5.64 9.96 ;
        RECT  4.56 4.08 5.64 4.56 ;
        RECT  4.56 3.00 5.04 4.56 ;
        RECT  2.28 2.94 2.88 3.54 ;
        RECT  1.26 11.58 1.86 12.18 ;
        RECT  1.32 10.44 1.80 12.18 ;
        LAYER via ;
        RECT  5.88 11.70 6.24 12.06 ;
        RECT  5.76 3.06 6.12 3.42 ;
        RECT  2.40 3.06 2.76 3.42 ;
        RECT  1.38 11.70 1.74 12.06 ;
        LAYER metal2 ;
        RECT  5.76 11.58 6.36 12.18 ;
        RECT  1.26 11.58 1.86 12.18 ;
        RECT  1.26 11.64 6.36 12.12 ;
        RECT  5.64 2.94 6.24 3.54 ;
        RECT  2.28 2.94 2.88 3.54 ;
        RECT  2.28 3.00 6.24 3.48 ;
    END
END lrp_1

MACRO lrp_2
    CLASS CORE ;
    FOREIGN lrp_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.04 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN rb
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal2 ;
        RECT  1.86 8.34 2.46 8.94 ;
        RECT  1.86 8.40 10.02 8.88 ;
        RECT  9.42 8.34 10.02 8.94 ;
        LAYER metal1 ;
        RECT  1.86 8.34 2.46 8.94 ;
        RECT  9.42 8.34 10.02 8.94 ;
        LAYER via ;
        RECT  1.98 8.46 2.34 8.82 ;
        RECT  9.54 8.46 9.90 8.82 ;
        END
    END rb
    PIN q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.40 6.24 13.20 6.72 ;
        RECT  12.72 5.16 13.20 7.80 ;
        RECT  12.96 2.76 13.44 5.64 ;
        RECT  12.96 7.32 13.44 12.36 ;
        END
    END q
    PIN ip
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 6.24 1.32 6.72 ;
        END
    END ip
    PIN ck
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER metal2 ;
        RECT  4.02 6.18 4.62 6.78 ;
        RECT  4.02 6.24 7.86 6.72 ;
        RECT  7.26 6.18 7.86 6.78 ;
        LAYER metal1 ;
        RECT  4.08 6.18 4.56 7.80 ;
        RECT  4.02 6.18 4.62 6.78 ;
        RECT  7.26 6.18 7.86 6.78 ;
        LAYER via ;
        RECT  4.14 6.30 4.50 6.66 ;
        RECT  7.38 6.30 7.74 6.66 ;
        END
    END ck
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.60 0.00 1.08 3.48 ;
        RECT  3.54 0.00 4.02 3.48 ;
        RECT  8.94 0.00 9.42 3.48 ;
        RECT  11.94 0.00 12.42 4.44 ;
        RECT  0.00 0.00 14.04 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.30 10.44 0.78 15.12 ;
        RECT  2.28 10.44 2.76 15.12 ;
        RECT  3.36 10.44 3.84 15.12 ;
        RECT  8.88 10.38 9.36 15.12 ;
        RECT  11.94 9.00 12.42 15.12 ;
        RECT  0.00 13.80 14.04 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  6.84 8.40 7.32 12.12 ;
        RECT  6.24 8.40 7.32 8.88 ;
        RECT  6.24 5.16 6.72 8.88 ;
        RECT  6.24 7.32 12.12 7.80 ;
        RECT  6.72 3.00 7.20 5.64 ;
        RECT  7.74 4.08 11.34 4.56 ;
        RECT  10.86 3.00 11.34 4.56 ;
        RECT  7.74 3.00 8.22 4.56 ;
        RECT  9.96 9.48 10.44 12.12 ;
        RECT  7.86 9.48 8.34 12.12 ;
        RECT  7.86 9.48 10.44 9.96 ;
        RECT  5.76 11.58 6.36 12.18 ;
        RECT  5.82 10.44 6.30 12.18 ;
        RECT  5.64 2.94 6.24 3.54 ;
        RECT  4.44 8.40 4.92 12.12 ;
        RECT  4.44 8.40 5.64 8.88 ;
        RECT  5.16 4.08 5.64 8.88 ;
        RECT  4.56 4.08 5.64 4.56 ;
        RECT  4.56 3.00 5.04 4.56 ;
        RECT  2.34 2.94 2.94 3.54 ;
        RECT  1.26 11.58 1.86 12.18 ;
        RECT  1.32 10.44 1.80 12.18 ;
        LAYER via ;
        RECT  5.88 11.70 6.24 12.06 ;
        RECT  5.76 3.06 6.12 3.42 ;
        RECT  2.46 3.06 2.82 3.42 ;
        RECT  1.38 11.70 1.74 12.06 ;
        LAYER metal2 ;
        RECT  5.76 11.58 6.36 12.18 ;
        RECT  1.26 11.58 1.86 12.18 ;
        RECT  1.26 11.64 6.36 12.12 ;
        RECT  5.64 2.94 6.24 3.54 ;
        RECT  2.34 2.94 2.94 3.54 ;
        RECT  2.34 3.00 6.24 3.48 ;
    END
END lrp_2

MACRO lrp_4
    CLASS CORE ;
    FOREIGN lrp_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.12 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN rb
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal2 ;
        RECT  1.86 8.34 2.46 8.94 ;
        RECT  1.86 8.40 10.02 8.88 ;
        RECT  9.42 8.34 10.02 8.94 ;
        LAYER metal1 ;
        RECT  1.86 8.34 2.46 8.94 ;
        RECT  9.42 8.34 10.02 8.94 ;
        LAYER via ;
        RECT  1.98 8.46 2.34 8.82 ;
        RECT  9.54 8.46 9.90 8.82 ;
        END
    END rb
    PIN q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.40 6.24 13.20 6.72 ;
        RECT  12.72 5.16 13.20 7.80 ;
        RECT  12.96 2.76 13.44 5.64 ;
        RECT  12.96 7.32 13.44 12.36 ;
        END
    END q
    PIN ip
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 6.24 1.32 6.72 ;
        END
    END ip
    PIN ck
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER metal2 ;
        RECT  4.02 6.18 4.62 6.78 ;
        RECT  4.02 6.24 7.86 6.72 ;
        RECT  7.26 6.18 7.86 6.78 ;
        LAYER metal1 ;
        RECT  4.08 6.18 4.56 7.80 ;
        RECT  4.02 6.18 4.62 6.78 ;
        RECT  7.26 6.18 7.86 6.78 ;
        LAYER via ;
        RECT  4.14 6.30 4.50 6.66 ;
        RECT  7.38 6.30 7.74 6.66 ;
        END
    END ck
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.60 0.00 1.08 3.48 ;
        RECT  3.54 0.00 4.02 3.48 ;
        RECT  8.94 0.00 9.42 3.48 ;
        RECT  11.94 0.00 12.42 4.44 ;
        RECT  13.98 0.00 14.46 4.44 ;
        RECT  0.00 0.00 15.12 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.30 10.20 0.78 15.12 ;
        RECT  2.28 10.20 2.76 15.12 ;
        RECT  3.36 10.20 3.84 15.12 ;
        RECT  8.88 10.32 9.36 15.12 ;
        RECT  11.94 9.00 12.42 15.12 ;
        RECT  13.98 9.00 14.46 15.12 ;
        RECT  0.00 13.80 15.12 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  6.84 8.40 7.32 12.36 ;
        RECT  6.24 8.40 7.32 8.88 ;
        RECT  6.24 5.16 6.72 8.88 ;
        RECT  6.24 7.32 12.12 7.80 ;
        RECT  6.72 3.06 7.20 5.64 ;
        RECT  7.74 4.08 11.34 4.56 ;
        RECT  10.86 3.06 11.34 4.56 ;
        RECT  7.74 3.06 8.22 4.56 ;
        RECT  9.96 9.48 10.44 12.36 ;
        RECT  7.86 9.48 8.34 12.36 ;
        RECT  7.86 9.48 10.44 9.96 ;
        RECT  5.82 10.20 6.30 12.36 ;
        RECT  5.76 11.58 6.36 12.18 ;
        RECT  5.64 2.94 6.24 3.54 ;
        RECT  4.44 8.40 4.92 12.36 ;
        RECT  4.44 8.40 5.64 8.88 ;
        RECT  5.16 4.08 5.64 8.88 ;
        RECT  4.56 4.08 5.64 4.56 ;
        RECT  4.56 3.00 5.04 4.56 ;
        RECT  2.28 2.94 2.88 3.54 ;
        RECT  1.32 10.20 1.80 12.36 ;
        RECT  1.26 11.58 1.86 12.18 ;
        LAYER via ;
        RECT  5.88 11.70 6.24 12.06 ;
        RECT  5.76 3.06 6.12 3.42 ;
        RECT  2.40 3.06 2.76 3.42 ;
        RECT  1.38 11.70 1.74 12.06 ;
        LAYER metal2 ;
        RECT  5.76 11.58 6.36 12.18 ;
        RECT  1.26 11.58 1.86 12.18 ;
        RECT  1.26 11.64 6.36 12.12 ;
        RECT  5.64 2.94 6.24 3.54 ;
        RECT  2.28 2.94 2.88 3.54 ;
        RECT  2.28 3.00 6.24 3.48 ;
    END
END lrp_4

MACRO lrsp_1
    CLASS CORE ;
    FOREIGN lrsp_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.20 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN s
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal2 ;
        RECT  1.86 5.10 2.46 5.70 ;
        RECT  1.86 5.16 10.02 5.64 ;
        RECT  9.42 5.10 10.02 5.70 ;
        LAYER metal1 ;
        RECT  1.86 5.10 2.46 5.70 ;
        RECT  9.42 5.10 10.02 5.70 ;
        LAYER via ;
        RECT  1.98 5.22 2.34 5.58 ;
        RECT  9.54 5.22 9.90 5.58 ;
        END
    END s
    PIN rb
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal2 ;
        RECT  2.94 9.42 3.54 10.02 ;
        RECT  2.94 9.48 12.18 9.96 ;
        RECT  11.58 9.42 12.18 10.02 ;
        LAYER metal1 ;
        RECT  2.94 9.42 3.54 10.02 ;
        RECT  11.58 9.42 12.18 10.02 ;
        LAYER via ;
        RECT  3.06 9.54 3.42 9.90 ;
        RECT  11.70 9.54 12.06 9.90 ;
        END
    END rb
    PIN q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.56 6.24 15.36 6.72 ;
        RECT  14.88 4.08 15.36 9.96 ;
        RECT  15.06 3.00 15.54 4.56 ;
        RECT  15.06 9.48 15.54 12.12 ;
        END
    END q
    PIN ip
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 6.24 1.32 6.72 ;
        END
    END ip
    PIN ck
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER metal2 ;
        RECT  5.10 8.34 5.70 8.94 ;
        RECT  5.10 8.40 8.94 8.88 ;
        RECT  8.34 8.34 8.94 8.94 ;
        LAYER metal1 ;
        RECT  5.10 8.34 5.70 8.94 ;
        RECT  8.34 8.34 8.94 8.94 ;
        LAYER via ;
        RECT  5.22 8.46 5.58 8.82 ;
        RECT  8.46 8.46 8.82 8.82 ;
        END
    END ck
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.38 0.00 1.86 3.48 ;
        RECT  4.62 0.00 5.10 3.48 ;
        RECT  10.92 0.00 11.40 3.48 ;
        RECT  14.04 0.00 14.52 3.48 ;
        RECT  0.00 0.00 16.20 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.66 10.44 1.14 15.12 ;
        RECT  3.36 10.44 3.84 15.12 ;
        RECT  4.44 10.44 4.92 15.12 ;
        RECT  10.80 10.44 11.28 15.12 ;
        RECT  14.04 10.44 14.52 15.12 ;
        RECT  0.00 13.80 16.20 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  7.92 9.48 8.40 12.12 ;
        RECT  7.32 9.48 8.40 9.96 ;
        RECT  7.32 5.10 7.80 9.96 ;
        RECT  7.32 7.32 14.28 7.80 ;
        RECT  7.80 3.00 8.28 5.58 ;
        RECT  12.84 2.94 13.44 3.54 ;
        RECT  9.96 4.08 12.36 4.56 ;
        RECT  11.88 3.00 12.36 4.56 ;
        RECT  9.96 3.00 10.44 4.56 ;
        RECT  11.76 11.58 12.36 12.18 ;
        RECT  11.82 10.44 12.30 12.18 ;
        RECT  8.88 11.58 9.48 12.18 ;
        RECT  8.94 10.44 9.42 12.18 ;
        RECT  8.76 2.94 9.36 3.54 ;
        RECT  6.84 11.58 7.44 12.18 ;
        RECT  6.90 10.44 7.38 12.18 ;
        RECT  6.72 2.94 7.32 3.54 ;
        RECT  5.52 9.48 6.00 12.12 ;
        RECT  5.52 9.48 6.72 9.96 ;
        RECT  6.24 4.08 6.72 9.96 ;
        RECT  5.64 4.08 6.72 4.56 ;
        RECT  5.64 3.00 6.12 4.56 ;
        RECT  3.36 2.94 3.96 3.54 ;
        RECT  2.34 11.58 2.94 12.18 ;
        RECT  2.40 10.44 2.88 12.18 ;
        RECT  0.42 4.08 2.82 4.56 ;
        RECT  2.34 3.00 2.82 4.56 ;
        RECT  0.42 3.00 0.90 4.56 ;
        LAYER via ;
        RECT  12.96 3.06 13.32 3.42 ;
        RECT  11.88 11.70 12.24 12.06 ;
        RECT  9.00 11.70 9.36 12.06 ;
        RECT  8.88 3.06 9.24 3.42 ;
        RECT  6.96 11.70 7.32 12.06 ;
        RECT  6.84 3.06 7.20 3.42 ;
        RECT  3.48 3.06 3.84 3.42 ;
        RECT  2.46 11.70 2.82 12.06 ;
        LAYER metal2 ;
        RECT  12.84 2.94 13.44 3.54 ;
        RECT  8.76 2.94 9.36 3.54 ;
        RECT  8.76 3.00 13.44 3.48 ;
        RECT  11.76 11.58 12.36 12.18 ;
        RECT  8.88 11.58 9.48 12.18 ;
        RECT  8.82 11.64 12.36 12.12 ;
        RECT  6.84 11.58 7.44 12.18 ;
        RECT  2.34 11.58 2.94 12.18 ;
        RECT  2.34 11.64 7.44 12.12 ;
        RECT  6.72 2.94 7.32 3.54 ;
        RECT  3.36 2.94 3.96 3.54 ;
        RECT  3.36 3.00 7.32 3.48 ;
    END
END lrsp_1

MACRO lrsp_2
    CLASS CORE ;
    FOREIGN lrsp_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.20 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN s
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal2 ;
        RECT  1.86 5.10 2.46 5.70 ;
        RECT  1.86 5.16 10.02 5.64 ;
        RECT  9.42 5.10 10.02 5.70 ;
        LAYER metal1 ;
        RECT  1.86 5.10 2.46 5.70 ;
        RECT  9.42 5.10 10.02 5.70 ;
        LAYER via ;
        RECT  1.98 5.22 2.34 5.58 ;
        RECT  9.54 5.22 9.90 5.58 ;
        END
    END s
    PIN rb
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal2 ;
        RECT  2.94 8.34 3.54 8.94 ;
        RECT  2.94 8.40 12.18 8.88 ;
        RECT  11.58 8.34 12.18 8.94 ;
        LAYER metal1 ;
        RECT  2.94 8.34 3.54 8.94 ;
        RECT  11.58 8.34 12.18 8.94 ;
        LAYER via ;
        RECT  3.06 8.46 3.42 8.82 ;
        RECT  11.70 8.46 12.06 8.82 ;
        END
    END rb
    PIN q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.56 6.24 15.36 6.72 ;
        RECT  14.88 4.50 15.36 8.70 ;
        RECT  15.06 2.76 15.54 4.98 ;
        RECT  15.06 8.22 15.54 12.36 ;
        END
    END q
    PIN ip
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 6.24 1.32 6.72 ;
        END
    END ip
    PIN ck
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER metal2 ;
        RECT  5.10 6.18 5.70 6.78 ;
        RECT  5.10 6.24 8.94 6.72 ;
        RECT  8.34 6.18 8.94 6.78 ;
        LAYER metal1 ;
        RECT  5.10 6.18 5.70 6.78 ;
        RECT  8.34 6.18 8.94 6.78 ;
        LAYER via ;
        RECT  5.22 6.30 5.58 6.66 ;
        RECT  8.46 6.30 8.82 6.66 ;
        END
    END ck
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.38 0.00 1.86 3.48 ;
        RECT  4.62 0.00 5.10 3.48 ;
        RECT  10.92 0.00 11.40 3.48 ;
        RECT  14.04 0.00 14.52 4.44 ;
        RECT  0.00 0.00 16.20 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.66 10.44 1.14 15.12 ;
        RECT  3.36 10.44 3.84 15.12 ;
        RECT  4.44 10.44 4.92 15.12 ;
        RECT  10.80 10.44 11.28 15.12 ;
        RECT  14.04 9.00 14.52 15.12 ;
        RECT  0.00 13.80 16.20 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  7.92 9.00 8.40 12.12 ;
        RECT  7.32 9.00 8.40 9.48 ;
        RECT  7.32 5.10 7.80 9.48 ;
        RECT  7.32 7.32 14.28 7.80 ;
        RECT  7.80 3.00 8.28 5.58 ;
        RECT  12.84 2.94 13.44 3.54 ;
        RECT  9.96 4.08 12.36 4.56 ;
        RECT  11.88 3.00 12.36 4.56 ;
        RECT  9.96 3.00 10.44 4.56 ;
        RECT  11.76 11.58 12.36 12.18 ;
        RECT  11.82 10.44 12.30 12.18 ;
        RECT  8.88 11.58 9.48 12.18 ;
        RECT  8.94 10.44 9.42 12.18 ;
        RECT  8.76 2.94 9.36 3.54 ;
        RECT  6.84 11.58 7.44 12.18 ;
        RECT  6.90 10.44 7.38 12.18 ;
        RECT  6.72 2.94 7.32 3.54 ;
        RECT  5.52 9.00 6.00 12.12 ;
        RECT  5.52 9.00 6.72 9.48 ;
        RECT  6.24 4.08 6.72 9.48 ;
        RECT  5.64 4.08 6.72 4.56 ;
        RECT  5.64 3.00 6.12 4.56 ;
        RECT  3.36 2.94 3.96 3.54 ;
        RECT  2.34 11.58 2.94 12.18 ;
        RECT  2.40 10.44 2.88 12.18 ;
        RECT  0.42 4.08 2.82 4.56 ;
        RECT  2.34 3.00 2.82 4.56 ;
        RECT  0.42 3.00 0.90 4.56 ;
        LAYER via ;
        RECT  12.96 3.06 13.32 3.42 ;
        RECT  11.88 11.70 12.24 12.06 ;
        RECT  9.00 11.70 9.36 12.06 ;
        RECT  8.88 3.06 9.24 3.42 ;
        RECT  6.96 11.70 7.32 12.06 ;
        RECT  6.84 3.06 7.20 3.42 ;
        RECT  3.48 3.06 3.84 3.42 ;
        RECT  2.46 11.70 2.82 12.06 ;
        LAYER metal2 ;
        RECT  12.84 2.94 13.44 3.54 ;
        RECT  8.76 2.94 9.36 3.54 ;
        RECT  8.76 3.00 13.44 3.48 ;
        RECT  11.76 11.58 12.36 12.18 ;
        RECT  8.88 11.58 9.48 12.18 ;
        RECT  8.82 11.64 12.36 12.12 ;
        RECT  6.84 11.58 7.44 12.18 ;
        RECT  2.34 11.58 2.94 12.18 ;
        RECT  2.34 11.64 7.44 12.12 ;
        RECT  6.72 2.94 7.32 3.54 ;
        RECT  3.36 2.94 3.96 3.54 ;
        RECT  3.36 3.00 7.32 3.48 ;
    END
END lrsp_2

MACRO lrsp_4
    CLASS CORE ;
    FOREIGN lrsp_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 17.28 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN s
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal2 ;
        RECT  1.86 5.10 2.46 5.70 ;
        RECT  1.86 5.16 10.02 5.64 ;
        RECT  9.42 5.10 10.02 5.70 ;
        LAYER metal1 ;
        RECT  1.86 5.10 2.46 5.70 ;
        RECT  9.42 5.10 10.02 5.70 ;
        LAYER via ;
        RECT  1.98 5.22 2.34 5.58 ;
        RECT  9.54 5.22 9.90 5.58 ;
        END
    END s
    PIN rb
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal2 ;
        RECT  2.94 8.34 3.54 8.94 ;
        RECT  2.94 8.40 12.18 8.88 ;
        RECT  11.58 8.34 12.18 8.94 ;
        LAYER metal1 ;
        RECT  2.94 8.34 3.54 8.94 ;
        RECT  11.58 8.34 12.18 8.94 ;
        LAYER via ;
        RECT  3.06 8.46 3.42 8.82 ;
        RECT  11.70 8.46 12.06 8.82 ;
        END
    END rb
    PIN q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.56 6.24 15.36 6.72 ;
        RECT  14.88 4.50 15.36 8.70 ;
        RECT  15.06 2.76 15.54 4.98 ;
        RECT  15.06 8.22 15.54 12.36 ;
        END
    END q
    PIN ip
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 6.24 1.32 6.72 ;
        END
    END ip
    PIN ck
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER metal2 ;
        RECT  5.10 6.18 5.70 6.78 ;
        RECT  5.10 6.24 8.94 6.72 ;
        RECT  8.34 6.18 8.94 6.78 ;
        LAYER metal1 ;
        RECT  5.10 6.18 5.70 6.78 ;
        RECT  8.34 6.18 8.94 6.78 ;
        LAYER via ;
        RECT  5.22 6.30 5.58 6.66 ;
        RECT  8.46 6.30 8.82 6.66 ;
        END
    END ck
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.38 0.00 1.86 3.54 ;
        RECT  4.62 0.00 5.10 3.54 ;
        RECT  10.92 0.00 11.40 3.54 ;
        RECT  14.04 0.00 14.52 4.44 ;
        RECT  16.08 0.00 16.56 4.44 ;
        RECT  0.00 0.00 17.28 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.66 9.96 1.14 15.12 ;
        RECT  3.36 9.96 3.84 15.12 ;
        RECT  4.44 9.96 4.92 15.12 ;
        RECT  10.80 9.96 11.28 15.12 ;
        RECT  14.04 9.00 14.52 15.12 ;
        RECT  16.08 9.00 16.56 15.12 ;
        RECT  0.00 13.80 17.28 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  7.92 9.00 8.40 12.12 ;
        RECT  7.32 9.00 8.40 9.48 ;
        RECT  7.32 5.10 7.80 9.48 ;
        RECT  7.32 7.32 14.28 7.80 ;
        RECT  7.80 3.06 8.28 5.58 ;
        RECT  12.84 2.94 13.44 3.54 ;
        RECT  9.96 4.08 12.36 4.56 ;
        RECT  11.88 3.06 12.36 4.56 ;
        RECT  9.96 3.06 10.44 4.56 ;
        RECT  11.76 11.58 12.36 12.18 ;
        RECT  11.82 9.96 12.30 12.18 ;
        RECT  8.88 11.58 9.48 12.18 ;
        RECT  8.94 9.96 9.42 12.18 ;
        RECT  8.76 2.94 9.36 3.54 ;
        RECT  6.84 11.58 7.44 12.18 ;
        RECT  6.90 9.96 7.38 12.18 ;
        RECT  6.72 2.94 7.32 3.54 ;
        RECT  5.52 9.00 6.00 12.12 ;
        RECT  5.52 9.00 6.72 9.48 ;
        RECT  6.24 4.08 6.72 9.48 ;
        RECT  5.64 4.08 6.72 4.56 ;
        RECT  5.64 3.06 6.12 4.56 ;
        RECT  3.36 2.94 3.96 3.54 ;
        RECT  2.34 11.58 2.94 12.18 ;
        RECT  2.40 9.96 2.88 12.18 ;
        RECT  0.42 4.08 2.82 4.56 ;
        RECT  2.34 3.06 2.82 4.56 ;
        RECT  0.42 3.06 0.90 4.56 ;
        LAYER via ;
        RECT  12.96 3.06 13.32 3.42 ;
        RECT  11.88 11.70 12.24 12.06 ;
        RECT  9.00 11.70 9.36 12.06 ;
        RECT  8.88 3.06 9.24 3.42 ;
        RECT  6.96 11.70 7.32 12.06 ;
        RECT  6.84 3.06 7.20 3.42 ;
        RECT  3.48 3.06 3.84 3.42 ;
        RECT  2.46 11.70 2.82 12.06 ;
        LAYER metal2 ;
        RECT  12.84 2.94 13.44 3.54 ;
        RECT  8.76 2.94 9.36 3.54 ;
        RECT  8.76 3.00 13.44 3.48 ;
        RECT  11.76 11.58 12.36 12.18 ;
        RECT  8.88 11.58 9.48 12.18 ;
        RECT  8.82 11.64 12.36 12.12 ;
        RECT  6.84 11.58 7.44 12.18 ;
        RECT  2.34 11.58 2.94 12.18 ;
        RECT  2.34 11.64 7.44 12.12 ;
        RECT  6.72 2.94 7.32 3.54 ;
        RECT  3.36 2.94 3.96 3.54 ;
        RECT  3.36 3.00 7.32 3.48 ;
    END
END lrsp_4

MACRO mux2_1
    CLASS CORE ;
    FOREIGN mux2_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.56 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN s
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal2 ;
        RECT  0.78 8.34 1.38 8.94 ;
        RECT  0.78 8.40 5.70 8.88 ;
        RECT  5.10 8.34 5.70 8.94 ;
        LAYER metal1 ;
        RECT  0.78 8.34 1.38 8.94 ;
        RECT  5.10 8.34 5.70 8.94 ;
        LAYER via ;
        RECT  0.90 8.46 1.26 8.82 ;
        RECT  5.22 8.46 5.58 8.82 ;
        END
    END s
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.24 4.08 6.72 9.96 ;
        RECT  6.60 3.00 7.08 5.04 ;
        RECT  6.60 9.00 7.08 12.36 ;
        END
    END op
    PIN ip2
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  3.00 6.24 3.48 6.72 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  5.16 7.32 5.64 7.80 ;
        END
    END ip1
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.26 0.00 1.74 3.48 ;
        RECT  4.68 0.00 5.16 3.48 ;
        RECT  5.64 0.00 6.12 3.48 ;
        RECT  0.00 0.00 7.56 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.26 10.68 1.74 15.12 ;
        RECT  4.68 10.68 5.16 15.12 ;
        RECT  5.64 10.68 6.12 15.12 ;
        RECT  0.00 13.80 7.56 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  5.10 5.10 5.70 5.70 ;
        RECT  3.00 7.32 3.48 12.36 ;
        RECT  3.00 7.32 4.56 7.80 ;
        RECT  4.08 4.32 4.56 7.80 ;
        RECT  4.08 6.24 5.64 6.72 ;
        RECT  2.94 4.32 4.56 4.80 ;
        RECT  2.94 3.00 3.42 4.80 ;
        RECT  0.30 9.48 0.78 12.36 ;
        RECT  0.30 9.48 2.40 9.96 ;
        RECT  1.92 7.32 2.40 9.96 ;
        RECT  0.84 7.32 2.40 7.80 ;
        RECT  0.84 5.16 1.32 7.80 ;
        RECT  1.86 5.10 2.46 5.70 ;
        RECT  0.30 5.16 2.46 5.64 ;
        RECT  0.30 3.00 0.78 5.64 ;
        LAYER via ;
        RECT  5.22 5.22 5.58 5.58 ;
        RECT  1.98 5.22 2.34 5.58 ;
        LAYER metal2 ;
        RECT  5.10 5.10 5.70 5.70 ;
        RECT  1.86 5.10 2.46 5.70 ;
        RECT  1.86 5.16 5.70 5.64 ;
    END
END mux2_1

MACRO mux2_2
    CLASS CORE ;
    FOREIGN mux2_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.56 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN s
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal2 ;
        RECT  0.78 8.34 1.38 8.94 ;
        RECT  0.78 8.40 5.70 8.88 ;
        RECT  5.10 8.34 5.70 8.94 ;
        LAYER metal1 ;
        RECT  0.78 8.34 1.38 8.94 ;
        RECT  5.10 8.34 5.70 8.94 ;
        LAYER via ;
        RECT  0.90 8.46 1.26 8.82 ;
        RECT  5.22 8.46 5.58 8.82 ;
        END
    END s
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.24 5.16 6.72 8.88 ;
        RECT  6.24 8.40 7.26 8.88 ;
        RECT  6.78 2.76 7.26 5.64 ;
        RECT  6.24 5.16 7.26 5.64 ;
        RECT  6.78 8.40 7.26 12.36 ;
        END
    END op
    PIN ip2
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  3.00 6.24 3.48 6.72 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  5.16 7.32 5.64 7.80 ;
        END
    END ip1
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.26 0.00 1.74 3.48 ;
        RECT  4.68 0.00 5.16 3.48 ;
        RECT  5.82 0.00 6.30 4.44 ;
        RECT  0.00 0.00 7.56 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.26 10.20 1.74 15.12 ;
        RECT  4.68 10.20 5.16 15.12 ;
        RECT  5.82 9.30 6.30 15.12 ;
        RECT  0.00 13.80 7.56 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  5.10 5.10 5.70 5.70 ;
        RECT  3.00 7.32 3.48 11.88 ;
        RECT  3.00 7.32 4.56 7.80 ;
        RECT  4.08 4.32 4.56 7.80 ;
        RECT  4.08 6.24 5.64 6.72 ;
        RECT  2.94 4.32 4.56 4.80 ;
        RECT  2.94 3.00 3.42 4.80 ;
        RECT  0.30 9.36 0.78 11.88 ;
        RECT  0.30 9.36 2.40 9.84 ;
        RECT  1.92 7.32 2.40 9.84 ;
        RECT  0.78 7.32 2.40 7.80 ;
        RECT  0.78 4.08 1.26 7.80 ;
        RECT  1.86 5.10 2.46 5.70 ;
        RECT  0.78 5.16 2.46 5.64 ;
        RECT  0.30 3.00 0.78 4.56 ;
        LAYER via ;
        RECT  5.22 5.22 5.58 5.58 ;
        RECT  1.98 5.22 2.34 5.58 ;
        LAYER metal2 ;
        RECT  5.10 5.10 5.70 5.70 ;
        RECT  1.86 5.10 2.46 5.70 ;
        RECT  1.86 5.16 5.70 5.64 ;
    END
END mux2_2

MACRO mux2_4
    CLASS CORE ;
    FOREIGN mux2_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.64 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN s
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal2 ;
        RECT  0.78 8.34 1.38 8.94 ;
        RECT  0.78 8.40 5.70 8.88 ;
        RECT  5.10 8.34 5.70 8.94 ;
        LAYER metal1 ;
        RECT  0.78 8.34 1.38 8.94 ;
        RECT  5.10 8.34 5.70 8.94 ;
        LAYER via ;
        RECT  0.90 8.46 1.26 8.82 ;
        RECT  5.22 8.46 5.58 8.82 ;
        END
    END s
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.90 2.76 7.38 5.64 ;
        RECT  6.90 8.40 7.38 12.36 ;
        RECT  7.32 5.16 7.80 8.88 ;
        END
    END op
    PIN ip2
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  3.00 6.24 3.48 6.72 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  5.16 7.32 5.64 7.80 ;
        END
    END ip1
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.26 0.00 1.74 3.48 ;
        RECT  4.68 0.00 5.16 3.48 ;
        RECT  5.94 0.00 6.42 4.44 ;
        RECT  7.86 0.00 8.34 4.44 ;
        RECT  0.00 0.00 8.64 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.26 10.50 1.74 15.12 ;
        RECT  4.68 10.50 5.16 15.12 ;
        RECT  5.94 9.30 6.42 15.12 ;
        RECT  7.86 9.30 8.34 15.12 ;
        RECT  0.00 13.80 8.64 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  3.00 7.32 3.48 12.12 ;
        RECT  3.00 7.32 4.56 7.80 ;
        RECT  4.08 4.32 4.56 7.80 ;
        RECT  4.08 6.24 6.72 6.72 ;
        RECT  2.94 4.32 4.56 4.80 ;
        RECT  2.94 3.00 3.42 4.80 ;
        RECT  5.10 5.10 5.70 5.70 ;
        RECT  0.30 9.36 0.78 12.12 ;
        RECT  0.30 9.36 2.40 9.84 ;
        RECT  1.92 7.32 2.40 9.84 ;
        RECT  0.84 7.32 2.40 7.80 ;
        RECT  0.84 5.16 1.32 7.80 ;
        RECT  1.86 5.10 2.46 5.70 ;
        RECT  0.30 5.16 2.46 5.64 ;
        RECT  0.30 3.00 0.78 5.64 ;
        LAYER via ;
        RECT  5.22 5.22 5.58 5.58 ;
        RECT  1.98 5.22 2.34 5.58 ;
        LAYER metal2 ;
        RECT  5.10 5.10 5.70 5.70 ;
        RECT  1.86 5.10 2.46 5.70 ;
        RECT  1.86 5.16 5.70 5.64 ;
    END
END mux2_4

MACRO mux3_2
    CLASS CORE ;
    FOREIGN mux3_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 19.44 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN s1
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal2 ;
        RECT  9.48 6.18 10.08 6.78 ;
        RECT  9.48 6.24 14.40 6.72 ;
        RECT  13.80 6.18 14.40 6.78 ;
        LAYER metal1 ;
        RECT  9.48 6.18 10.08 6.78 ;
        RECT  13.80 6.18 14.40 6.78 ;
        LAYER via ;
        RECT  9.60 6.30 9.96 6.66 ;
        RECT  13.92 6.30 14.28 6.66 ;
        END
    END s1
    PIN s0
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal2 ;
        RECT  1.92 7.26 2.52 7.86 ;
        RECT  1.92 7.32 6.84 7.80 ;
        RECT  6.24 7.26 6.84 7.86 ;
        LAYER metal1 ;
        RECT  1.92 7.26 2.52 7.86 ;
        RECT  6.24 7.26 6.84 7.86 ;
        LAYER via ;
        RECT  2.04 7.38 2.40 7.74 ;
        RECT  6.36 7.38 6.72 7.74 ;
        END
    END s0
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  17.64 2.76 18.12 5.64 ;
        RECT  17.64 8.40 18.12 12.36 ;
        RECT  17.64 5.16 18.66 5.64 ;
        RECT  18.18 5.16 18.66 8.88 ;
        RECT  17.64 8.40 18.66 8.88 ;
        END
    END op
    PIN ip3
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  16.02 5.16 16.50 5.64 ;
        END
    END ip3
    PIN ip2
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  8.46 7.32 8.94 7.80 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.90 6.24 1.38 6.72 ;
        END
    END ip1
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.44 0.00 1.92 4.44 ;
        RECT  9.00 0.00 9.48 4.44 ;
        RECT  16.56 0.00 17.04 4.44 ;
        RECT  0.00 0.00 19.44 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.44 9.00 1.92 15.12 ;
        RECT  9.00 9.00 9.48 15.12 ;
        RECT  16.56 9.00 17.04 15.12 ;
        RECT  0.00 13.80 19.44 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  17.04 7.26 17.64 7.86 ;
        RECT  15.48 9.00 15.96 12.36 ;
        RECT  13.86 7.32 14.34 12.36 ;
        RECT  13.86 11.70 15.96 12.18 ;
        RECT  13.80 8.34 14.40 8.94 ;
        RECT  13.86 7.32 15.42 7.80 ;
        RECT  14.94 5.16 15.42 7.80 ;
        RECT  13.86 5.16 15.42 5.64 ;
        RECT  13.86 2.76 14.34 5.64 ;
        RECT  15.48 2.76 15.96 4.44 ;
        RECT  13.86 2.94 15.96 3.42 ;
        RECT  12.78 2.76 13.26 12.36 ;
        RECT  12.72 7.26 13.32 7.86 ;
        RECT  11.70 2.76 12.18 12.36 ;
        RECT  11.64 8.34 12.24 8.94 ;
        RECT  10.08 8.40 10.56 12.36 ;
        RECT  10.08 8.40 11.10 8.88 ;
        RECT  10.62 5.16 11.10 8.88 ;
        RECT  10.08 5.16 11.10 5.64 ;
        RECT  10.08 2.76 10.56 5.64 ;
        RECT  7.92 8.40 8.40 12.36 ;
        RECT  6.18 8.40 6.66 12.36 ;
        RECT  6.18 8.40 8.40 8.88 ;
        RECT  7.38 5.16 7.86 8.88 ;
        RECT  6.18 6.24 7.86 6.72 ;
        RECT  6.18 2.76 6.66 6.72 ;
        RECT  7.38 5.16 8.40 5.64 ;
        RECT  7.92 2.76 8.40 5.64 ;
        RECT  5.10 2.76 5.58 12.36 ;
        RECT  5.04 8.34 5.64 8.94 ;
        RECT  4.02 2.76 4.50 12.36 ;
        RECT  3.96 11.58 4.56 12.18 ;
        RECT  3.96 2.94 4.56 3.54 ;
        RECT  2.52 8.40 3.00 12.36 ;
        RECT  2.52 8.40 3.54 8.88 ;
        RECT  3.06 5.16 3.54 8.88 ;
        RECT  2.52 5.16 3.54 5.64 ;
        RECT  2.52 2.76 3.00 5.64 ;
        RECT  0.36 2.76 0.84 4.44 ;
        RECT  0.30 2.94 0.90 3.54 ;
        RECT  0.36 9.00 0.84 12.36 ;
        RECT  0.30 11.58 0.90 12.18 ;
        LAYER via ;
        RECT  17.16 7.38 17.52 7.74 ;
        RECT  13.92 8.46 14.28 8.82 ;
        RECT  12.84 7.38 13.20 7.74 ;
        RECT  11.76 8.46 12.12 8.82 ;
        RECT  5.16 8.46 5.52 8.82 ;
        RECT  4.08 3.06 4.44 3.42 ;
        RECT  4.08 11.70 4.44 12.06 ;
        RECT  0.42 3.06 0.78 3.42 ;
        RECT  0.42 11.70 0.78 12.06 ;
        LAYER metal2 ;
        RECT  17.04 7.26 17.64 7.86 ;
        RECT  12.72 7.26 13.32 7.86 ;
        RECT  12.72 7.32 17.64 7.80 ;
        RECT  13.80 8.34 14.40 8.94 ;
        RECT  11.64 8.34 12.24 8.94 ;
        RECT  5.04 8.34 5.64 8.94 ;
        RECT  5.04 8.40 12.24 8.88 ;
        RECT  3.96 2.94 4.56 3.54 ;
        RECT  0.30 2.94 0.90 3.54 ;
        RECT  0.30 3.00 4.56 3.48 ;
        RECT  3.96 11.58 4.56 12.18 ;
        RECT  0.30 11.58 0.90 12.18 ;
        RECT  0.30 11.64 4.56 12.12 ;
    END
END mux3_2

MACRO mux4_2
    CLASS CORE ;
    FOREIGN mux4_2 0.06 0 ;
    ORIGIN -0.06 0.00 ;
    SIZE 24.84 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN s1
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal2 ;
        RECT  9.48 6.18 10.08 6.78 ;
        RECT  9.48 6.24 14.40 6.72 ;
        RECT  13.80 6.18 14.40 6.78 ;
        LAYER metal1 ;
        RECT  9.48 6.18 10.08 6.78 ;
        RECT  13.80 6.18 14.40 6.78 ;
        LAYER via ;
        RECT  9.60 6.30 9.96 6.66 ;
        RECT  13.92 6.30 14.28 6.66 ;
        END
    END s1
    PIN s0
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal2 ;
        RECT  1.92 7.26 2.52 7.86 ;
        RECT  6.24 7.26 6.84 7.86 ;
        RECT  18.12 7.26 18.72 7.86 ;
        RECT  1.92 7.32 20.88 7.80 ;
        RECT  20.28 7.26 20.88 7.86 ;
        LAYER metal1 ;
        RECT  1.92 7.26 2.52 7.86 ;
        RECT  6.24 7.26 6.84 7.86 ;
        RECT  18.12 7.26 18.72 7.86 ;
        RECT  20.28 7.26 20.88 7.86 ;
        LAYER via ;
        RECT  2.04 7.38 2.40 7.74 ;
        RECT  6.36 7.38 6.72 7.74 ;
        RECT  18.24 7.38 18.60 7.74 ;
        RECT  20.40 7.38 20.76 7.74 ;
        END
    END s0
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  23.58 2.76 24.06 12.36 ;
        END
    END op
    PIN ip4
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  21.42 5.16 21.90 5.64 ;
        END
    END ip4
    PIN ip3
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  16.02 6.24 16.50 6.72 ;
        END
    END ip3
    PIN ip2
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  8.46 6.24 8.94 6.72 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.90 6.24 1.38 6.72 ;
        END
    END ip1
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.44 0.00 1.92 4.44 ;
        RECT  9.00 0.00 9.48 4.44 ;
        RECT  15.48 0.00 15.96 4.44 ;
        RECT  22.50 0.00 22.98 4.44 ;
        RECT  0.06 0.00 24.90 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.44 9.00 1.92 15.12 ;
        RECT  9.00 9.00 9.48 15.12 ;
        RECT  15.48 9.00 15.96 15.12 ;
        RECT  22.50 9.00 22.98 15.12 ;
        RECT  0.06 13.80 24.90 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  22.44 7.26 23.04 7.86 ;
        RECT  21.42 6.24 21.90 12.36 ;
        RECT  19.80 10.68 20.28 12.36 ;
        RECT  19.80 11.70 21.90 12.18 ;
        RECT  20.34 6.24 21.90 6.72 ;
        RECT  20.34 2.76 20.82 6.72 ;
        RECT  21.42 2.76 21.90 4.44 ;
        RECT  20.34 2.94 21.90 3.42 ;
        RECT  18.72 8.34 19.20 12.36 ;
        RECT  18.66 8.34 19.26 8.94 ;
        RECT  19.26 2.76 19.74 8.88 ;
        RECT  18.12 5.10 18.72 5.70 ;
        RECT  17.64 10.68 18.12 12.36 ;
        RECT  16.56 8.40 17.04 12.36 ;
        RECT  16.56 11.70 18.12 12.18 ;
        RECT  16.56 8.40 17.58 8.88 ;
        RECT  17.10 5.16 17.58 8.88 ;
        RECT  16.56 5.16 17.58 5.64 ;
        RECT  16.56 2.76 17.04 5.64 ;
        RECT  18.18 2.76 18.66 3.60 ;
        RECT  16.56 2.94 18.66 3.42 ;
        RECT  13.86 7.32 14.34 12.36 ;
        RECT  13.80 8.34 14.40 8.94 ;
        RECT  13.86 7.32 15.42 7.80 ;
        RECT  14.94 5.16 15.42 7.80 ;
        RECT  13.86 5.16 15.42 5.64 ;
        RECT  13.86 2.76 14.34 5.64 ;
        RECT  12.78 2.76 13.26 12.36 ;
        RECT  12.72 9.42 13.32 10.02 ;
        RECT  11.70 2.76 12.18 12.36 ;
        RECT  11.64 8.34 12.24 8.94 ;
        RECT  10.08 8.40 10.56 12.36 ;
        RECT  10.08 8.40 11.10 8.88 ;
        RECT  10.62 5.16 11.10 8.88 ;
        RECT  10.08 5.16 11.10 5.64 ;
        RECT  10.08 2.76 10.56 5.64 ;
        RECT  7.92 8.40 8.40 12.36 ;
        RECT  6.18 8.40 6.66 12.36 ;
        RECT  6.18 8.40 8.40 8.88 ;
        RECT  7.38 5.16 7.86 8.88 ;
        RECT  6.18 5.16 8.40 5.64 ;
        RECT  7.92 2.76 8.40 5.64 ;
        RECT  6.18 2.76 6.66 5.64 ;
        RECT  5.10 2.76 5.58 12.36 ;
        RECT  5.04 8.34 5.64 8.94 ;
        RECT  4.02 2.76 4.50 12.36 ;
        RECT  3.96 11.58 4.56 12.18 ;
        RECT  3.96 2.94 4.56 3.54 ;
        RECT  2.52 8.40 3.00 12.36 ;
        RECT  2.52 8.40 3.54 8.88 ;
        RECT  3.06 5.10 3.54 8.88 ;
        RECT  3.00 5.10 3.60 5.70 ;
        RECT  2.52 2.76 3.00 5.64 ;
        RECT  0.36 2.76 0.84 4.44 ;
        RECT  0.30 2.94 0.90 3.54 ;
        RECT  0.36 9.00 0.84 12.36 ;
        RECT  0.30 11.58 0.90 12.18 ;
        LAYER via ;
        RECT  22.56 7.38 22.92 7.74 ;
        RECT  18.78 8.46 19.14 8.82 ;
        RECT  18.24 5.22 18.60 5.58 ;
        RECT  13.92 8.46 14.28 8.82 ;
        RECT  12.84 9.54 13.20 9.90 ;
        RECT  11.76 8.46 12.12 8.82 ;
        RECT  5.16 8.46 5.52 8.82 ;
        RECT  4.08 3.06 4.44 3.42 ;
        RECT  4.08 11.70 4.44 12.06 ;
        RECT  3.12 5.22 3.48 5.58 ;
        RECT  0.42 3.06 0.78 3.42 ;
        RECT  0.42 11.70 0.78 12.06 ;
        LAYER metal2 ;
        RECT  12.72 9.42 13.32 10.02 ;
        RECT  12.72 9.48 22.98 9.96 ;
        RECT  22.50 7.26 22.98 9.96 ;
        RECT  22.44 7.26 23.04 7.86 ;
        RECT  18.66 8.34 19.26 8.94 ;
        RECT  13.80 8.34 14.40 8.94 ;
        RECT  13.80 8.40 19.26 8.88 ;
        RECT  18.12 5.10 18.72 5.70 ;
        RECT  3.00 5.10 3.60 5.70 ;
        RECT  3.00 5.16 18.72 5.64 ;
        RECT  11.64 8.34 12.24 8.94 ;
        RECT  5.04 8.34 5.64 8.94 ;
        RECT  5.04 8.40 12.24 8.88 ;
        RECT  3.96 2.94 4.56 3.54 ;
        RECT  0.30 2.94 0.90 3.54 ;
        RECT  0.30 3.00 4.56 3.48 ;
        RECT  3.96 11.58 4.56 12.18 ;
        RECT  0.30 11.58 0.90 12.18 ;
        RECT  0.30 11.64 4.56 12.12 ;
    END
END mux4_2

MACRO nand2_1
    CLASS CORE ;
    FOREIGN nand2_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.32 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.86 9.48 2.34 12.24 ;
        RECT  3.00 3.00 3.48 9.96 ;
        RECT  1.86 9.48 3.48 9.96 ;
        END
    END op
    PIN ip2
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  1.92 6.24 2.40 6.72 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 7.32 1.32 7.80 ;
        END
    END ip1
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.26 0.00 1.74 3.48 ;
        RECT  0.00 0.00 4.32 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.84 10.68 1.32 15.12 ;
        RECT  2.94 10.68 3.42 15.12 ;
        RECT  0.00 13.80 4.32 15.12 ;
        END
    END vdd
END nand2_1

MACRO nand2_2
    CLASS CORE ;
    FOREIGN nand2_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.32 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.92 8.40 2.40 12.30 ;
        RECT  3.00 2.88 3.48 8.88 ;
        RECT  1.92 8.40 3.48 8.88 ;
        END
    END op
    PIN ip2
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  1.92 6.24 2.40 6.72 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 7.32 1.32 7.80 ;
        END
    END ip1
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.32 0.00 1.80 4.44 ;
        RECT  0.00 0.00 4.32 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.90 9.00 1.38 15.12 ;
        RECT  3.00 9.48 3.48 15.12 ;
        RECT  0.00 13.80 4.32 15.12 ;
        END
    END vdd
END nand2_2

MACRO nand2_4
    CLASS CORE ;
    FOREIGN nand2_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.48 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.92 8.40 2.40 12.30 ;
        RECT  3.00 2.88 3.48 8.88 ;
        RECT  3.00 2.88 3.54 4.44 ;
        RECT  1.92 8.40 4.50 8.88 ;
        RECT  4.02 8.40 4.50 12.30 ;
        END
    END op
    PIN ip2
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  1.92 6.24 2.40 6.72 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal2 ;
        RECT  0.78 7.26 1.38 7.86 ;
        RECT  0.78 7.32 5.70 7.80 ;
        RECT  5.10 7.26 5.70 7.86 ;
        LAYER metal1 ;
        RECT  0.78 7.26 1.38 7.86 ;
        RECT  5.10 7.26 5.70 7.86 ;
        LAYER via ;
        RECT  0.90 7.38 1.26 7.74 ;
        RECT  5.22 7.38 5.58 7.74 ;
        END
    END ip1
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.32 0.00 1.80 4.44 ;
        RECT  4.86 0.00 5.34 4.44 ;
        RECT  0.00 0.00 6.48 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.90 9.42 1.38 15.12 ;
        RECT  3.00 9.48 3.48 15.12 ;
        RECT  5.10 9.48 5.58 15.12 ;
        RECT  0.00 13.80 6.48 15.12 ;
        END
    END vdd
END nand2_4

MACRO nand3_1
    CLASS CORE ;
    FOREIGN nand3_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.40 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.86 9.48 2.34 12.24 ;
        RECT  3.00 3.00 3.48 9.96 ;
        RECT  1.86 9.48 4.44 9.96 ;
        RECT  3.00 3.00 4.14 3.48 ;
        RECT  3.96 9.48 4.44 12.24 ;
        END
    END op
    PIN ip3
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  4.08 5.16 4.56 5.64 ;
        END
    END ip3
    PIN ip2
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  1.92 6.24 2.40 6.72 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 7.32 1.32 7.80 ;
        END
    END ip1
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.20 0.00 1.68 3.60 ;
        RECT  0.00 0.00 5.40 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.84 10.56 1.32 15.12 ;
        RECT  2.94 10.56 3.42 15.12 ;
        RECT  0.00 13.80 5.40 15.12 ;
        END
    END vdd
END nand3_1

MACRO nand3_2
    CLASS CORE ;
    FOREIGN nand3_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.40 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.84 8.40 1.32 12.30 ;
        RECT  1.92 7.32 2.40 8.88 ;
        RECT  0.84 8.40 3.42 8.88 ;
        RECT  2.94 8.40 3.42 12.30 ;
        RECT  3.00 4.08 3.48 7.80 ;
        RECT  1.92 7.32 3.48 7.80 ;
        RECT  3.66 2.82 4.14 4.56 ;
        RECT  3.00 4.08 4.14 4.56 ;
        END
    END op
    PIN ip3
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  4.08 5.16 4.56 5.64 ;
        END
    END ip3
    PIN ip2
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  1.92 6.24 2.40 6.72 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 7.32 1.32 7.80 ;
        END
    END ip1
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.20 0.00 1.68 4.44 ;
        RECT  0.00 0.00 5.40 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.86 9.48 2.34 15.12 ;
        RECT  3.96 9.12 4.44 15.12 ;
        RECT  0.00 13.80 5.40 15.12 ;
        END
    END vdd
END nand3_2

MACRO nand3_4
    CLASS CORE ;
    FOREIGN nand3_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.64 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.84 8.40 1.32 12.24 ;
        RECT  1.92 7.32 2.40 8.88 ;
        RECT  0.84 8.40 3.42 8.88 ;
        RECT  2.94 8.40 3.42 12.24 ;
        RECT  3.00 4.08 3.48 7.80 ;
        RECT  1.92 7.32 3.48 7.80 ;
        RECT  3.66 2.94 4.14 4.56 ;
        RECT  3.00 4.08 4.14 4.56 ;
        END
    END op
    PIN ip3
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  4.08 5.16 4.56 5.64 ;
        END
    END ip3
    PIN ip2
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal2 ;
        RECT  1.86 6.18 2.46 6.78 ;
        RECT  1.86 6.24 5.70 6.72 ;
        RECT  5.10 6.18 5.70 6.78 ;
        LAYER metal1 ;
        RECT  1.86 6.18 2.46 6.78 ;
        RECT  5.10 6.18 5.70 6.78 ;
        LAYER via ;
        RECT  1.98 6.30 2.34 6.66 ;
        RECT  5.22 6.30 5.58 6.66 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal2 ;
        RECT  0.78 7.26 1.38 7.86 ;
        RECT  0.78 7.32 7.86 7.80 ;
        RECT  7.26 7.26 7.86 7.86 ;
        LAYER metal1 ;
        RECT  0.78 7.26 1.38 7.86 ;
        RECT  7.26 7.26 7.86 7.86 ;
        LAYER via ;
        RECT  0.90 7.38 1.26 7.74 ;
        RECT  7.38 7.38 7.74 7.74 ;
        END
    END ip1
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.20 0.00 1.68 4.44 ;
        RECT  6.12 0.00 6.60 4.44 ;
        RECT  0.00 0.00 8.64 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.86 9.48 2.34 15.12 ;
        RECT  3.96 9.48 4.44 15.12 ;
        RECT  6.06 9.48 6.54 15.12 ;
        RECT  0.00 13.80 8.64 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  7.08 8.40 7.56 12.24 ;
        RECT  4.98 8.40 5.46 12.24 ;
        RECT  4.98 8.40 7.56 8.88 ;
    END
END nand3_4

MACRO nand4_1
    CLASS CORE ;
    FOREIGN nand4_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.40 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.32 9.54 1.80 12.18 ;
        RECT  3.00 7.32 3.48 10.02 ;
        RECT  1.32 9.54 4.02 10.02 ;
        RECT  3.54 9.54 4.02 12.18 ;
        RECT  4.08 2.88 4.56 7.80 ;
        RECT  3.00 7.32 4.56 7.80 ;
        RECT  4.08 2.88 4.68 3.72 ;
        END
    END op
    PIN ip4
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  4.08 8.40 4.56 8.88 ;
        END
    END ip4
    PIN ip3
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  3.00 6.24 3.48 6.72 ;
        END
    END ip3
    PIN ip2
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  1.92 8.40 2.40 8.88 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 5.16 1.32 5.64 ;
        END
    END ip1
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.96 0.00 1.44 3.60 ;
        RECT  0.00 0.00 5.40 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.30 10.50 0.78 15.12 ;
        RECT  2.40 10.50 2.88 15.12 ;
        RECT  4.62 10.50 5.10 15.12 ;
        RECT  0.00 13.80 5.40 15.12 ;
        END
    END vdd
END nand4_1

MACRO nand4_2
    CLASS CORE ;
    FOREIGN nand4_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.40 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.32 8.40 1.80 12.30 ;
        RECT  3.00 6.24 3.48 8.88 ;
        RECT  1.32 8.40 4.02 8.88 ;
        RECT  3.54 8.40 4.02 12.30 ;
        RECT  4.08 2.76 4.56 6.72 ;
        RECT  3.00 6.24 4.56 6.72 ;
        RECT  4.08 2.76 4.68 4.20 ;
        END
    END op
    PIN ip4
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  4.08 7.32 4.56 7.80 ;
        END
    END ip4
    PIN ip3
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  3.00 5.16 3.48 5.64 ;
        END
    END ip3
    PIN ip2
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  1.92 7.32 2.40 7.80 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 5.16 1.32 5.64 ;
        END
    END ip1
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.96 0.00 1.44 4.08 ;
        RECT  0.00 0.00 5.40 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.30 9.42 0.78 15.12 ;
        RECT  2.40 9.48 2.88 15.12 ;
        RECT  4.62 9.42 5.10 15.12 ;
        RECT  0.00 13.80 5.40 15.12 ;
        END
    END vdd
END nand4_2

MACRO nand4_4
    CLASS CORE ;
    FOREIGN nand4_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.80 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.04 2.76 8.52 5.64 ;
        RECT  8.04 8.40 8.52 12.24 ;
        RECT  8.40 5.16 8.88 8.88 ;
        END
    END op
    PIN ip4
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  4.08 6.24 4.56 6.72 ;
        END
    END ip4
    PIN ip3
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  3.00 5.16 3.48 5.64 ;
        END
    END ip3
    PIN ip2
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  1.92 5.16 2.40 5.64 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 7.32 1.32 7.80 ;
        END
    END ip1
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  4.20 0.00 4.68 4.08 ;
        RECT  6.84 0.00 7.32 4.08 ;
        RECT  9.36 0.00 9.84 4.08 ;
        RECT  0.00 0.00 10.80 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.30 9.42 0.78 15.12 ;
        RECT  2.40 9.48 2.88 15.12 ;
        RECT  4.62 9.42 5.10 15.12 ;
        RECT  6.84 9.42 7.32 15.12 ;
        RECT  9.30 9.42 9.78 15.12 ;
        RECT  0.00 13.80 10.80 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  5.76 8.40 6.24 12.24 ;
        RECT  6.24 6.24 6.72 8.88 ;
        RECT  6.24 7.32 7.80 7.80 ;
        RECT  5.34 6.24 6.72 6.72 ;
        RECT  5.34 2.76 5.82 6.72 ;
        RECT  3.54 8.40 4.02 12.30 ;
        RECT  1.32 8.40 1.80 12.30 ;
        RECT  1.32 8.40 4.02 8.88 ;
        RECT  2.94 6.24 3.42 8.88 ;
        RECT  2.94 7.32 5.64 7.80 ;
        RECT  0.96 6.24 3.42 6.72 ;
        RECT  0.96 2.82 1.44 6.72 ;
    END
END nand4_4

MACRO nor2_1
    CLASS CORE ;
    FOREIGN nor2_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 3.24 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.84 7.32 1.32 9.96 ;
        RECT  1.38 3.00 1.86 5.64 ;
        RECT  1.38 5.16 2.40 5.64 ;
        RECT  1.92 5.16 2.40 7.80 ;
        RECT  0.84 7.32 2.40 7.80 ;
        RECT  0.84 9.48 2.94 9.96 ;
        RECT  2.46 9.48 2.94 12.30 ;
        END
    END op
    PIN ip2
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  1.92 8.40 2.40 8.88 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 6.24 1.32 6.72 ;
        END
    END ip1
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.30 0.00 0.78 3.60 ;
        RECT  2.46 0.00 2.94 3.60 ;
        RECT  0.00 0.00 3.24 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.66 10.62 1.14 15.12 ;
        RECT  0.00 13.80 3.24 15.12 ;
        END
    END vdd
END nor2_1

MACRO nor2_2
    CLASS CORE ;
    FOREIGN nor2_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 3.24 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.84 6.24 1.32 8.88 ;
        RECT  1.44 2.76 1.92 4.56 ;
        RECT  1.92 4.08 2.40 6.72 ;
        RECT  0.84 6.24 2.40 6.72 ;
        RECT  0.84 8.40 2.94 8.88 ;
        RECT  2.46 8.40 2.94 12.24 ;
        END
    END op
    PIN ip2
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  1.92 7.32 2.40 7.80 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 5.16 1.32 5.64 ;
        END
    END ip1
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.42 0.00 0.90 3.66 ;
        RECT  2.46 0.00 2.94 3.60 ;
        RECT  0.00 0.00 3.24 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.72 9.24 1.20 15.12 ;
        RECT  0.00 13.80 3.24 15.12 ;
        END
    END vdd
END nor2_2

MACRO nor2_4
    CLASS CORE ;
    FOREIGN nor2_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.56 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.92 2.88 2.40 5.64 ;
        RECT  3.00 5.16 3.48 12.24 ;
        RECT  5.22 2.88 5.70 5.64 ;
        RECT  1.92 5.16 6.72 5.64 ;
        RECT  6.24 5.16 6.72 12.24 ;
        END
    END op
    PIN ip2
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal2 ;
        RECT  1.86 7.26 2.46 7.86 ;
        RECT  1.86 7.32 5.70 7.80 ;
        RECT  5.10 7.26 5.70 7.86 ;
        LAYER metal1 ;
        RECT  1.86 7.26 2.46 7.86 ;
        RECT  5.10 7.26 5.70 7.86 ;
        LAYER via ;
        RECT  1.98 7.38 2.34 7.74 ;
        RECT  5.22 7.38 5.58 7.74 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal2 ;
        RECT  0.78 6.18 1.38 6.78 ;
        RECT  0.78 6.24 4.62 6.72 ;
        RECT  4.02 6.18 4.62 6.78 ;
        LAYER metal1 ;
        RECT  0.78 6.18 1.38 6.78 ;
        RECT  4.02 6.18 4.62 6.78 ;
        LAYER via ;
        RECT  0.90 6.30 1.26 6.66 ;
        RECT  4.14 6.30 4.50 6.66 ;
        END
    END ip1
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.84 0.00 1.32 4.26 ;
        RECT  3.00 0.00 3.48 4.26 ;
        RECT  4.14 0.00 4.62 4.26 ;
        RECT  6.24 0.00 6.72 4.26 ;
        RECT  0.00 0.00 7.56 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.20 9.24 1.68 15.12 ;
        RECT  4.44 9.24 4.92 15.12 ;
        RECT  0.00 13.80 7.56 15.12 ;
        END
    END vdd
END nor2_4

MACRO nor3_1
    CLASS CORE ;
    FOREIGN nor3_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.32 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.50 3.00 1.98 4.56 ;
        RECT  1.92 4.08 2.40 6.72 ;
        RECT  1.92 6.24 3.48 6.72 ;
        RECT  3.00 6.24 3.48 12.06 ;
        RECT  3.00 10.38 3.60 12.06 ;
        RECT  3.54 3.00 4.02 4.56 ;
        RECT  1.50 4.08 4.02 4.56 ;
        END
    END op
    PIN ip3
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  3.00 5.16 3.48 5.64 ;
        END
    END ip3
    PIN ip2
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  1.92 7.32 2.40 7.80 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 6.24 1.32 6.72 ;
        END
    END ip1
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.48 0.00 0.96 3.60 ;
        RECT  2.58 0.00 3.06 3.60 ;
        RECT  0.00 0.00 4.32 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.72 10.38 1.20 15.12 ;
        RECT  0.00 13.80 4.32 15.12 ;
        END
    END vdd
END nor3_1

MACRO nor3_2
    CLASS CORE ;
    FOREIGN nor3_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.32 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.32 2.76 1.80 4.56 ;
        RECT  1.92 4.08 2.40 6.72 ;
        RECT  1.92 6.24 3.48 6.72 ;
        RECT  3.00 6.24 3.48 8.88 ;
        RECT  3.24 2.76 3.72 4.56 ;
        RECT  1.32 4.08 3.72 4.56 ;
        RECT  3.24 8.40 3.72 12.36 ;
        END
    END op
    PIN ip3
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  3.00 5.16 3.48 5.64 ;
        END
    END ip3
    PIN ip2
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  1.92 7.32 2.40 7.80 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 6.24 1.32 6.72 ;
        END
    END ip1
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.36 0.00 0.84 4.08 ;
        RECT  2.28 0.00 2.76 3.72 ;
        RECT  0.00 0.00 4.32 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.72 9.00 1.20 15.12 ;
        RECT  0.00 13.80 4.32 15.12 ;
        END
    END vdd
END nor3_2

MACRO nor3_4
    CLASS CORE ;
    FOREIGN nor3_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.56 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.44 3.00 1.92 5.64 ;
        RECT  3.00 5.16 3.48 8.88 ;
        RECT  3.48 8.40 3.96 12.36 ;
        RECT  3.60 3.00 4.08 5.64 ;
        RECT  5.70 3.00 6.18 5.64 ;
        RECT  1.44 5.16 6.18 5.64 ;
        END
    END op
    PIN ip3
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  4.08 6.24 4.56 6.72 ;
        END
    END ip3
    PIN ip2
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal2 ;
        RECT  1.86 7.26 2.46 7.86 ;
        RECT  1.86 7.32 5.70 7.80 ;
        RECT  5.10 7.26 5.70 7.86 ;
        LAYER metal1 ;
        RECT  1.86 7.26 2.46 7.86 ;
        RECT  5.10 7.26 5.70 7.86 ;
        LAYER via ;
        RECT  1.98 7.38 2.34 7.74 ;
        RECT  5.22 7.38 5.58 7.74 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal2 ;
        RECT  0.78 8.34 1.38 8.94 ;
        RECT  0.78 8.40 6.78 8.88 ;
        RECT  6.18 8.34 6.78 8.94 ;
        LAYER metal1 ;
        RECT  0.78 8.34 1.38 8.94 ;
        RECT  6.18 8.34 6.78 8.94 ;
        LAYER via ;
        RECT  0.90 8.46 1.26 8.82 ;
        RECT  6.30 8.46 6.66 8.82 ;
        END
    END ip1
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.36 0.00 0.84 4.44 ;
        RECT  2.58 0.00 3.06 4.44 ;
        RECT  4.62 0.00 5.10 4.44 ;
        RECT  6.78 0.00 7.26 4.44 ;
        RECT  0.00 0.00 7.56 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.02 9.30 1.50 15.12 ;
        RECT  6.00 9.30 6.48 15.12 ;
        RECT  0.00 13.80 7.56 15.12 ;
        END
    END vdd
END nor3_4

MACRO nor4_1
    CLASS CORE ;
    FOREIGN nor4_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.40 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.38 3.00 1.86 4.56 ;
        RECT  3.00 4.08 3.48 6.72 ;
        RECT  3.54 3.00 4.02 4.56 ;
        RECT  1.38 4.08 4.02 4.56 ;
        RECT  3.00 6.24 4.56 6.72 ;
        RECT  4.08 6.24 4.56 11.70 ;
        RECT  3.84 10.38 4.56 11.70 ;
        END
    END op
    PIN ip4
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  4.08 5.16 4.56 5.64 ;
        END
    END ip4
    PIN ip3
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  3.00 7.32 3.48 7.80 ;
        END
    END ip3
    PIN ip2
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  1.92 6.24 2.40 6.72 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 8.40 1.32 8.88 ;
        END
    END ip1
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.30 0.00 0.78 3.60 ;
        RECT  2.46 0.00 2.94 3.60 ;
        RECT  4.62 0.00 5.10 3.60 ;
        RECT  0.00 0.00 5.40 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.66 10.44 1.14 15.12 ;
        RECT  0.00 13.80 5.40 15.12 ;
        END
    END vdd
END nor4_1

MACRO nor4_2
    CLASS CORE ;
    FOREIGN nor4_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.40 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal2 ;
        RECT  1.32 2.94 1.92 3.54 ;
        RECT  1.32 3.06 4.08 3.42 ;
        RECT  3.48 2.94 4.08 3.54 ;
        LAYER metal1 ;
        RECT  3.54 2.88 4.02 4.44 ;
        RECT  3.48 2.94 4.08 3.54 ;
        RECT  1.38 2.94 1.86 5.64 ;
        RECT  1.32 2.94 1.92 3.54 ;
        RECT  1.38 5.16 3.48 5.64 ;
        RECT  3.00 5.16 3.48 6.72 ;
        RECT  3.00 6.24 4.56 6.72 ;
        RECT  4.08 6.24 4.56 12.36 ;
        RECT  3.84 9.06 4.56 12.36 ;
        LAYER via ;
        RECT  1.44 3.06 1.80 3.42 ;
        RECT  3.60 3.06 3.96 3.42 ;
        END
    END op
    PIN ip4
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  4.08 5.16 4.56 5.64 ;
        END
    END ip4
    PIN ip3
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  3.00 7.32 3.48 7.80 ;
        END
    END ip3
    PIN ip2
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  1.92 6.24 2.40 6.72 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 7.32 1.32 7.80 ;
        END
    END ip1
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.30 0.00 0.78 4.44 ;
        RECT  2.46 0.00 2.94 4.44 ;
        RECT  4.62 0.00 5.10 4.44 ;
        RECT  0.00 0.00 5.40 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.66 9.00 1.14 15.12 ;
        RECT  0.00 13.80 5.40 15.12 ;
        END
    END vdd
END nor4_2

MACRO nor4_4
    CLASS CORE ;
    FOREIGN nor4_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.80 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.88 2.76 9.36 5.64 ;
        RECT  8.88 8.40 9.36 12.36 ;
        RECT  8.88 5.16 9.96 5.64 ;
        RECT  9.48 5.16 9.96 8.88 ;
        RECT  8.88 8.40 9.96 8.88 ;
        END
    END op
    PIN ip4
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  4.08 5.16 4.56 5.64 ;
        END
    END ip4
    PIN ip3
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  3.00 7.32 3.48 7.80 ;
        END
    END ip3
    PIN ip2
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  1.92 6.24 2.40 6.72 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 7.32 1.32 7.80 ;
        END
    END ip1
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.30 0.00 0.78 4.44 ;
        RECT  2.46 0.00 2.94 4.44 ;
        RECT  4.62 0.00 5.10 4.44 ;
        RECT  5.70 0.00 6.18 4.44 ;
        RECT  7.80 0.00 8.28 4.44 ;
        RECT  9.96 0.00 10.44 4.44 ;
        RECT  0.00 0.00 10.80 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.66 9.00 1.14 15.12 ;
        RECT  5.70 9.00 6.18 15.12 ;
        RECT  7.80 9.24 8.28 15.12 ;
        RECT  9.90 9.24 10.38 15.12 ;
        RECT  0.00 13.80 10.80 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  6.72 8.40 7.20 12.36 ;
        RECT  6.72 8.40 7.80 8.88 ;
        RECT  7.32 5.16 7.80 8.88 ;
        RECT  7.32 7.32 8.88 7.80 ;
        RECT  6.72 5.16 7.80 5.64 ;
        RECT  6.72 2.76 7.20 5.64 ;
        RECT  3.84 6.24 4.32 12.36 ;
        RECT  3.84 7.32 6.72 7.80 ;
        RECT  3.00 6.24 4.32 6.72 ;
        RECT  3.00 5.16 3.48 6.72 ;
        RECT  1.38 5.16 3.48 5.64 ;
        RECT  1.38 2.94 1.86 5.64 ;
        RECT  1.32 2.94 1.92 3.54 ;
        RECT  3.54 2.94 4.02 4.44 ;
        RECT  3.48 2.94 4.08 3.54 ;
        LAYER via ;
        RECT  3.60 3.06 3.96 3.42 ;
        RECT  1.44 3.06 1.80 3.42 ;
        LAYER metal2 ;
        RECT  3.48 2.94 4.08 3.54 ;
        RECT  1.32 2.94 1.92 3.54 ;
        RECT  1.32 3.06 4.08 3.42 ;
    END
END nor4_4

MACRO not_ab_or_c_or_d
    CLASS CORE ;
    FOREIGN not_ab_or_c_or_d 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.56 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.00 2.88 3.48 4.56 ;
        RECT  3.00 4.08 5.64 4.56 ;
        RECT  5.16 2.88 5.64 7.80 ;
        RECT  5.16 7.32 6.72 7.80 ;
        RECT  6.24 7.32 6.72 12.24 ;
        END
    END op
    PIN ip4
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  6.24 5.16 6.72 5.64 ;
        END
    END ip4
    PIN ip3
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  4.08 7.32 4.56 7.80 ;
        END
    END ip3
    PIN ip2
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  3.00 6.24 3.48 6.72 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 5.16 1.32 5.64 ;
        END
    END ip1
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.84 0.00 1.32 3.54 ;
        RECT  4.08 0.00 4.56 3.72 ;
        RECT  6.24 0.00 6.72 3.72 ;
        RECT  0.00 0.00 7.56 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.84 10.56 1.32 15.12 ;
        RECT  3.00 10.56 3.48 15.12 ;
        RECT  0.00 13.80 7.56 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  4.08 9.48 4.56 12.24 ;
        RECT  1.92 9.48 2.40 12.24 ;
        RECT  1.92 9.48 4.56 9.96 ;
    END
END not_ab_or_c_or_d

MACRO or2_1
    CLASS CORE ;
    FOREIGN or2_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.40 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.08 3.00 4.56 12.36 ;
        RECT  4.08 3.00 4.68 3.66 ;
        RECT  4.08 10.80 4.68 12.36 ;
        END
    END op
    PIN ip2
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  1.92 7.32 2.40 7.80 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 5.16 1.32 5.64 ;
        END
    END ip1
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.84 0.00 1.32 3.48 ;
        RECT  3.00 0.00 3.48 3.48 ;
        RECT  0.00 0.00 5.40 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  3.00 10.80 3.48 15.12 ;
        RECT  0.00 13.80 5.40 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  1.20 8.40 1.68 12.36 ;
        RECT  0.84 6.24 1.32 8.88 ;
        RECT  0.84 6.24 3.48 6.72 ;
        RECT  1.92 3.00 2.40 6.72 ;
    END
END or2_1

MACRO or2_2
    CLASS CORE ;
    FOREIGN or2_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.40 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.08 2.76 4.56 12.36 ;
        RECT  4.08 2.76 4.68 4.32 ;
        RECT  4.08 9.00 4.68 12.36 ;
        END
    END op
    PIN ip2
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  1.92 7.32 2.40 7.80 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 5.16 1.32 5.64 ;
        END
    END ip1
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.84 0.00 1.32 4.20 ;
        RECT  3.00 0.00 3.48 4.32 ;
        RECT  0.00 0.00 5.40 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  3.00 9.00 3.48 15.12 ;
        RECT  0.00 13.80 5.40 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  1.20 8.40 1.68 12.36 ;
        RECT  0.84 6.24 1.32 8.88 ;
        RECT  0.84 6.24 3.48 6.72 ;
        RECT  1.92 2.76 2.40 6.72 ;
    END
END or2_2

MACRO or2_4
    CLASS CORE ;
    FOREIGN or2_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.40 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.42 7.32 3.90 12.36 ;
        RECT  3.54 2.76 4.02 5.64 ;
        RECT  3.54 5.16 4.56 5.64 ;
        RECT  4.08 5.16 4.56 7.80 ;
        RECT  3.42 7.32 4.56 7.80 ;
        END
    END op
    PIN ip2
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  1.92 7.32 2.40 7.80 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 5.16 1.32 5.64 ;
        END
    END ip1
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.30 0.00 0.78 4.14 ;
        RECT  2.46 0.00 2.94 3.72 ;
        RECT  4.62 0.00 5.10 4.14 ;
        RECT  0.00 0.00 5.40 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.34 9.00 2.82 15.12 ;
        RECT  4.44 9.00 4.92 15.12 ;
        RECT  0.00 13.80 5.40 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  0.48 8.40 0.96 12.36 ;
        RECT  0.84 6.24 1.32 8.88 ;
        RECT  0.84 6.24 3.48 6.72 ;
        RECT  1.92 4.08 2.40 6.72 ;
        RECT  1.38 4.08 2.40 4.56 ;
        RECT  1.38 2.76 1.86 4.56 ;
    END
END or2_4

MACRO or3_1
    CLASS CORE ;
    FOREIGN or3_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.48 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.08 7.32 4.56 9.96 ;
        RECT  4.08 9.48 5.64 9.96 ;
        RECT  5.16 5.10 5.64 7.80 ;
        RECT  4.08 7.32 5.64 7.80 ;
        RECT  5.16 9.48 5.64 12.24 ;
        RECT  5.70 3.00 6.18 5.64 ;
        RECT  5.16 5.10 6.18 5.64 ;
        END
    END op
    PIN ip3
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  4.08 6.24 4.56 6.72 ;
        END
    END ip3
    PIN ip2
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  1.92 7.32 2.40 7.80 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 6.24 1.32 6.72 ;
        END
    END ip1
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.46 0.00 2.94 3.48 ;
        RECT  4.62 0.00 5.10 3.48 ;
        RECT  0.00 0.00 6.48 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  4.02 10.56 4.50 15.12 ;
        RECT  0.00 13.80 6.48 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  5.10 8.34 5.70 8.94 ;
        RECT  1.56 10.56 2.04 12.24 ;
        RECT  1.56 10.56 3.48 11.04 ;
        RECT  3.00 4.08 3.48 11.04 ;
        RECT  2.94 8.34 3.54 8.94 ;
        RECT  1.38 4.08 4.02 4.56 ;
        RECT  3.54 3.00 4.02 4.56 ;
        RECT  1.38 3.00 1.86 4.56 ;
        LAYER via ;
        RECT  5.22 8.46 5.58 8.82 ;
        RECT  3.06 8.46 3.42 8.82 ;
        LAYER metal2 ;
        RECT  5.10 8.34 5.70 8.94 ;
        RECT  2.94 8.34 3.54 8.94 ;
        RECT  2.94 8.40 5.70 8.88 ;
    END
END or3_1

MACRO or3_2
    CLASS CORE ;
    FOREIGN or3_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.48 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.08 6.24 4.56 8.88 ;
        RECT  4.08 8.40 5.64 8.88 ;
        RECT  5.16 8.40 5.64 12.36 ;
        RECT  5.70 2.76 6.18 6.72 ;
        RECT  4.08 6.24 6.18 6.72 ;
        END
    END op
    PIN ip3
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  4.08 5.16 4.56 5.64 ;
        END
    END ip3
    PIN ip2
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  1.92 6.24 2.40 6.72 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 7.32 1.32 7.80 ;
        END
    END ip1
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.46 0.00 2.94 3.72 ;
        RECT  4.62 0.00 5.10 4.08 ;
        RECT  0.00 0.00 6.48 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  4.02 9.24 4.50 15.12 ;
        RECT  0.00 13.80 6.48 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  5.10 7.26 5.70 7.86 ;
        RECT  1.56 8.40 2.04 12.36 ;
        RECT  1.56 8.40 3.48 8.88 ;
        RECT  3.00 4.08 3.48 8.88 ;
        RECT  2.94 7.26 3.54 7.86 ;
        RECT  1.38 4.08 4.02 4.56 ;
        RECT  3.54 2.76 4.02 4.56 ;
        RECT  1.38 2.76 1.86 4.56 ;
        LAYER via ;
        RECT  5.22 7.38 5.58 7.74 ;
        RECT  3.06 7.38 3.42 7.74 ;
        LAYER metal2 ;
        RECT  5.10 7.26 5.70 7.86 ;
        RECT  2.94 7.26 3.54 7.86 ;
        RECT  2.94 7.32 5.70 7.80 ;
    END
END or3_2

MACRO or3_4
    CLASS CORE ;
    FOREIGN or3_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.56 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.16 6.24 5.64 12.36 ;
        RECT  5.70 2.76 6.18 6.72 ;
        RECT  5.16 6.24 6.18 6.72 ;
        END
    END op
    PIN ip3
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  4.08 5.16 4.56 5.64 ;
        END
    END ip3
    PIN ip2
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  1.92 6.24 2.40 6.72 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 5.16 1.32 5.64 ;
        END
    END ip1
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.46 0.00 2.94 3.72 ;
        RECT  4.62 0.00 5.10 4.08 ;
        RECT  6.78 0.00 7.26 4.08 ;
        RECT  0.00 0.00 7.56 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  4.02 9.00 4.50 15.12 ;
        RECT  6.24 9.00 6.72 15.12 ;
        RECT  0.00 13.80 7.56 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  6.18 7.26 6.78 7.86 ;
        RECT  1.56 8.40 2.04 12.36 ;
        RECT  1.56 8.40 3.48 8.88 ;
        RECT  3.00 4.08 3.48 8.88 ;
        RECT  2.94 7.26 3.54 7.86 ;
        RECT  1.38 4.08 4.02 4.56 ;
        RECT  3.54 2.76 4.02 4.56 ;
        RECT  1.38 2.76 1.86 4.56 ;
        LAYER via ;
        RECT  6.30 7.38 6.66 7.74 ;
        RECT  3.06 7.38 3.42 7.74 ;
        LAYER metal2 ;
        RECT  6.18 7.26 6.78 7.86 ;
        RECT  2.94 7.26 3.54 7.86 ;
        RECT  2.94 7.32 6.78 7.80 ;
    END
END or3_4

MACRO or4_1
    CLASS CORE ;
    FOREIGN or4_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.48 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.08 7.32 4.56 10.86 ;
        RECT  4.08 10.38 5.52 10.86 ;
        RECT  5.04 10.38 5.52 12.36 ;
        RECT  5.16 4.08 5.64 7.80 ;
        RECT  4.08 7.32 5.64 7.80 ;
        RECT  5.70 3.00 6.18 4.56 ;
        RECT  5.16 4.08 6.18 4.56 ;
        END
    END op
    PIN ip4
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  4.08 5.16 4.56 5.64 ;
        END
    END ip4
    PIN ip3
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  3.00 7.32 3.48 7.80 ;
        END
    END ip3
    PIN ip2
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  1.92 5.16 2.40 5.64 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 8.40 1.32 8.88 ;
        END
    END ip1
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.30 0.00 0.78 3.48 ;
        RECT  2.46 0.00 2.94 3.48 ;
        RECT  4.62 0.00 5.10 3.42 ;
        RECT  0.00 0.00 6.48 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  3.90 11.22 4.38 15.12 ;
        RECT  0.00 13.80 6.48 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  5.10 9.42 5.70 10.02 ;
        RECT  0.72 9.48 1.20 12.36 ;
        RECT  1.86 9.42 2.46 10.02 ;
        RECT  0.72 9.48 2.46 9.96 ;
        RECT  1.92 6.24 2.40 10.02 ;
        RECT  1.92 6.24 3.48 6.72 ;
        RECT  3.00 4.08 3.48 6.72 ;
        RECT  1.38 4.08 4.02 4.56 ;
        RECT  3.54 3.00 4.02 4.56 ;
        RECT  1.38 3.00 1.86 4.56 ;
        LAYER via ;
        RECT  5.22 9.54 5.58 9.90 ;
        RECT  1.98 9.54 2.34 9.90 ;
        LAYER metal2 ;
        RECT  5.10 9.42 5.70 10.02 ;
        RECT  1.86 9.42 2.46 10.02 ;
        RECT  1.86 9.48 5.70 9.96 ;
    END
END or4_1

MACRO or4_2
    CLASS CORE ;
    FOREIGN or4_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.48 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.08 6.24 4.56 8.88 ;
        RECT  4.08 8.40 5.88 8.88 ;
        RECT  5.16 4.44 5.64 6.72 ;
        RECT  4.08 6.24 5.64 6.72 ;
        RECT  5.40 8.40 5.88 12.36 ;
        RECT  5.70 2.76 6.18 4.92 ;
        RECT  5.16 4.44 6.18 4.92 ;
        END
    END op
    PIN ip4
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  4.08 5.16 4.56 5.64 ;
        END
    END ip4
    PIN ip3
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  3.00 6.24 3.48 6.72 ;
        END
    END ip3
    PIN ip2
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  1.92 5.16 2.40 5.64 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 7.32 1.32 7.80 ;
        END
    END ip1
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.30 0.00 0.78 3.78 ;
        RECT  2.46 0.00 2.94 3.78 ;
        RECT  4.62 0.00 5.10 4.08 ;
        RECT  0.00 0.00 6.48 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  4.44 9.24 4.92 15.12 ;
        RECT  0.00 13.80 6.48 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  5.10 7.26 5.70 7.86 ;
        RECT  1.32 8.40 1.80 12.36 ;
        RECT  1.32 8.40 2.40 8.88 ;
        RECT  1.92 6.24 2.40 8.88 ;
        RECT  1.86 7.26 2.46 7.86 ;
        RECT  0.84 6.24 2.40 6.72 ;
        RECT  0.84 4.14 1.32 6.72 ;
        RECT  0.84 4.14 4.02 4.62 ;
        RECT  3.54 2.76 4.02 4.62 ;
        RECT  1.38 2.76 1.86 4.62 ;
        LAYER via ;
        RECT  5.22 7.38 5.58 7.74 ;
        RECT  1.98 7.38 2.34 7.74 ;
        LAYER metal2 ;
        RECT  5.10 7.26 5.70 7.86 ;
        RECT  1.86 7.26 2.46 7.86 ;
        RECT  1.86 7.32 5.70 7.80 ;
    END
END or4_2

MACRO or4_4
    CLASS CORE ;
    FOREIGN or4_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.56 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.40 8.40 5.88 12.36 ;
        RECT  5.70 2.76 6.18 4.92 ;
        RECT  5.70 4.44 6.72 4.92 ;
        RECT  6.24 4.44 6.72 8.88 ;
        RECT  5.40 8.40 6.72 8.88 ;
        END
    END op
    PIN ip4
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  4.08 5.16 4.56 5.64 ;
        END
    END ip4
    PIN ip3
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  3.00 6.24 3.48 6.72 ;
        END
    END ip3
    PIN ip2
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  1.92 5.16 2.40 5.64 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal1 ;
        RECT  0.84 7.32 1.32 7.80 ;
        END
    END ip1
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.30 0.00 0.78 3.78 ;
        RECT  2.46 0.00 2.94 3.78 ;
        RECT  4.62 0.00 5.10 4.14 ;
        RECT  6.66 0.00 7.14 4.08 ;
        RECT  0.00 0.00 7.56 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  4.44 9.00 4.92 15.12 ;
        RECT  6.42 9.24 6.90 15.12 ;
        RECT  0.00 13.80 7.56 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  5.10 7.26 5.70 7.86 ;
        RECT  1.32 8.40 1.80 12.36 ;
        RECT  1.32 8.40 2.40 8.88 ;
        RECT  1.92 6.24 2.40 8.88 ;
        RECT  1.86 7.26 2.46 7.86 ;
        RECT  0.84 6.24 2.40 6.72 ;
        RECT  0.84 4.14 1.32 6.72 ;
        RECT  0.84 4.14 4.02 4.62 ;
        RECT  3.54 2.76 4.02 4.62 ;
        RECT  1.38 2.76 1.86 4.62 ;
        LAYER via ;
        RECT  5.22 7.38 5.58 7.74 ;
        RECT  1.98 7.38 2.34 7.74 ;
        LAYER metal2 ;
        RECT  5.10 7.26 5.70 7.86 ;
        RECT  1.86 7.26 2.46 7.86 ;
        RECT  1.86 7.32 5.70 7.80 ;
    END
END or4_4

MACRO xnor2_1
    CLASS CORE ;
    FOREIGN xnor2_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.72 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.40 4.08 8.88 9.96 ;
        RECT  8.40 9.48 9.42 9.96 ;
        RECT  8.94 3.00 9.42 4.56 ;
        RECT  8.40 4.08 9.42 4.56 ;
        RECT  8.94 9.48 9.42 12.12 ;
        END
    END op
    PIN ip2
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal2 ;
        RECT  0.78 6.18 1.38 6.78 ;
        RECT  0.78 6.24 5.70 6.72 ;
        RECT  5.10 6.18 5.70 6.78 ;
        LAYER metal1 ;
        RECT  0.78 6.18 1.38 6.78 ;
        RECT  5.10 6.18 5.70 6.78 ;
        LAYER via ;
        RECT  0.90 6.30 1.26 6.66 ;
        RECT  5.22 6.30 5.58 6.66 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal2 ;
        RECT  2.94 8.34 3.54 8.94 ;
        RECT  2.94 8.40 7.86 8.88 ;
        RECT  7.26 8.34 7.86 8.94 ;
        LAYER metal1 ;
        RECT  2.94 8.34 3.54 8.94 ;
        RECT  7.26 8.34 7.86 8.94 ;
        LAYER via ;
        RECT  3.06 8.46 3.42 8.82 ;
        RECT  7.38 8.46 7.74 8.82 ;
        END
    END ip1
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.42 0.00 0.90 3.48 ;
        RECT  3.42 0.00 3.90 3.48 ;
        RECT  6.84 0.00 7.32 3.48 ;
        RECT  7.98 0.00 8.46 3.48 ;
        RECT  0.00 0.00 9.72 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.42 10.44 0.90 15.12 ;
        RECT  3.42 10.44 3.90 15.12 ;
        RECT  6.84 10.44 7.32 15.12 ;
        RECT  7.98 10.44 8.46 15.12 ;
        RECT  0.00 13.80 9.72 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  7.26 5.10 7.86 5.70 ;
        RECT  7.26 7.26 7.86 7.86 ;
        RECT  5.16 7.80 5.64 12.12 ;
        RECT  5.16 7.80 6.72 8.28 ;
        RECT  6.24 4.32 6.72 8.28 ;
        RECT  6.24 6.24 7.80 6.72 ;
        RECT  5.10 4.32 6.72 4.80 ;
        RECT  5.10 3.00 5.58 4.80 ;
        RECT  2.46 9.48 2.94 12.12 ;
        RECT  2.46 9.48 4.56 9.96 ;
        RECT  4.08 4.08 4.56 9.96 ;
        RECT  4.02 5.10 4.62 5.70 ;
        RECT  2.46 4.08 4.56 4.56 ;
        RECT  2.46 3.00 2.94 4.56 ;
        RECT  1.38 8.40 1.86 12.12 ;
        RECT  1.38 8.40 2.40 8.88 ;
        RECT  1.92 5.10 2.40 8.88 ;
        RECT  1.86 7.26 2.46 7.86 ;
        RECT  1.38 5.10 2.40 5.58 ;
        RECT  1.38 3.00 1.86 5.58 ;
        LAYER via ;
        RECT  7.38 5.22 7.74 5.58 ;
        RECT  7.38 7.38 7.74 7.74 ;
        RECT  4.14 5.22 4.50 5.58 ;
        RECT  1.98 7.38 2.34 7.74 ;
        LAYER metal2 ;
        RECT  7.26 5.10 7.86 5.70 ;
        RECT  4.02 5.10 4.62 5.70 ;
        RECT  4.02 5.16 7.86 5.64 ;
        RECT  7.26 7.26 7.86 7.86 ;
        RECT  1.86 7.26 2.46 7.86 ;
        RECT  1.86 7.32 7.86 7.80 ;
    END
END xnor2_1

MACRO xnor2_2
    CLASS CORE ;
    FOREIGN xnor2_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.72 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.40 5.16 8.88 8.88 ;
        RECT  8.40 8.40 9.42 8.88 ;
        RECT  8.94 2.76 9.42 5.64 ;
        RECT  8.40 5.16 9.42 5.64 ;
        RECT  8.94 8.40 9.42 12.36 ;
        END
    END op
    PIN ip2
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal2 ;
        RECT  0.78 6.18 1.38 6.78 ;
        RECT  0.78 6.24 5.70 6.72 ;
        RECT  5.10 6.18 5.70 6.78 ;
        LAYER metal1 ;
        RECT  0.78 6.18 1.38 6.78 ;
        RECT  5.10 6.18 5.70 6.78 ;
        LAYER via ;
        RECT  0.90 6.30 1.26 6.66 ;
        RECT  5.22 6.30 5.58 6.66 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal2 ;
        RECT  2.94 8.34 3.54 8.94 ;
        RECT  2.94 8.40 7.86 8.88 ;
        RECT  7.26 8.34 7.86 8.94 ;
        LAYER metal1 ;
        RECT  2.94 8.34 3.54 8.94 ;
        RECT  7.26 8.34 7.86 8.94 ;
        LAYER via ;
        RECT  3.06 8.46 3.42 8.82 ;
        RECT  7.38 8.46 7.74 8.82 ;
        END
    END ip1
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.42 0.00 0.90 3.48 ;
        RECT  3.42 0.00 3.90 3.48 ;
        RECT  6.84 0.00 7.32 3.48 ;
        RECT  7.98 0.00 8.46 4.44 ;
        RECT  0.00 0.00 9.72 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.42 10.38 0.90 15.12 ;
        RECT  3.42 10.38 3.90 15.12 ;
        RECT  6.84 10.38 7.32 15.12 ;
        RECT  7.98 9.30 8.46 15.12 ;
        RECT  0.00 13.80 9.72 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  7.26 5.10 7.86 5.70 ;
        RECT  7.26 7.26 7.86 7.86 ;
        RECT  5.16 7.80 5.64 12.06 ;
        RECT  5.16 7.80 6.72 8.28 ;
        RECT  6.24 4.32 6.72 8.28 ;
        RECT  6.24 6.24 7.80 6.72 ;
        RECT  5.10 4.32 6.72 4.80 ;
        RECT  5.10 3.00 5.58 4.80 ;
        RECT  2.46 9.48 2.94 12.06 ;
        RECT  2.46 9.48 4.56 9.96 ;
        RECT  4.08 4.08 4.56 9.96 ;
        RECT  4.02 5.10 4.62 5.70 ;
        RECT  2.46 4.08 4.56 4.56 ;
        RECT  2.46 3.00 2.94 4.56 ;
        RECT  1.38 8.40 1.86 12.06 ;
        RECT  1.38 8.40 2.40 8.88 ;
        RECT  1.92 5.10 2.40 8.88 ;
        RECT  1.86 7.26 2.46 7.86 ;
        RECT  1.38 5.10 2.40 5.58 ;
        RECT  1.38 3.00 1.86 5.58 ;
        LAYER via ;
        RECT  7.38 5.22 7.74 5.58 ;
        RECT  7.38 7.38 7.74 7.74 ;
        RECT  4.14 5.22 4.50 5.58 ;
        RECT  1.98 7.38 2.34 7.74 ;
        LAYER metal2 ;
        RECT  7.26 5.10 7.86 5.70 ;
        RECT  4.02 5.10 4.62 5.70 ;
        RECT  4.02 5.16 7.86 5.64 ;
        RECT  7.26 7.26 7.86 7.86 ;
        RECT  1.86 7.26 2.46 7.86 ;
        RECT  1.86 7.32 7.86 7.80 ;
    END
END xnor2_2

MACRO xor2_1
    CLASS CORE ;
    FOREIGN xor2_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.64 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.10 3.00 5.58 4.80 ;
        RECT  5.16 9.48 5.64 12.24 ;
        RECT  5.10 4.32 6.72 4.80 ;
        RECT  6.24 4.32 6.72 9.96 ;
        RECT  5.16 9.48 6.72 9.96 ;
        END
    END op
    PIN ip2
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal2 ;
        RECT  0.78 7.26 1.38 7.86 ;
        RECT  0.78 7.32 5.70 7.80 ;
        RECT  5.10 7.26 5.70 7.86 ;
        LAYER metal1 ;
        RECT  0.78 7.26 1.38 7.86 ;
        RECT  5.10 7.26 5.70 7.86 ;
        LAYER via ;
        RECT  0.90 7.38 1.26 7.74 ;
        RECT  5.22 7.38 5.58 7.74 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal2 ;
        RECT  2.94 8.34 3.54 8.94 ;
        RECT  2.94 8.40 7.86 8.88 ;
        RECT  7.26 8.34 7.86 8.94 ;
        LAYER metal1 ;
        RECT  2.94 8.34 3.54 8.94 ;
        RECT  7.26 8.34 7.86 8.94 ;
        LAYER via ;
        RECT  3.06 8.46 3.42 8.82 ;
        RECT  7.38 8.46 7.74 8.82 ;
        END
    END ip1
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.42 0.00 0.90 3.48 ;
        RECT  3.42 0.00 3.90 3.48 ;
        RECT  6.84 0.00 7.32 3.48 ;
        RECT  0.00 0.00 8.64 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.42 10.56 0.90 15.12 ;
        RECT  3.42 10.56 3.90 15.12 ;
        RECT  6.84 10.56 7.32 15.12 ;
        RECT  0.00 13.80 8.64 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  7.26 5.10 7.86 5.70 ;
        RECT  7.26 6.18 7.86 6.78 ;
        RECT  2.46 9.48 2.94 12.24 ;
        RECT  2.46 9.48 4.56 9.96 ;
        RECT  4.08 4.08 4.56 9.96 ;
        RECT  4.02 5.10 4.62 5.70 ;
        RECT  2.46 4.08 4.56 4.56 ;
        RECT  2.46 3.00 2.94 4.56 ;
        RECT  1.38 8.40 1.86 12.24 ;
        RECT  1.38 8.40 2.40 8.88 ;
        RECT  1.92 5.10 2.40 8.88 ;
        RECT  1.86 6.18 2.46 6.78 ;
        RECT  1.38 5.10 2.40 5.58 ;
        RECT  1.38 3.00 1.86 5.58 ;
        LAYER via ;
        RECT  7.38 5.22 7.74 5.58 ;
        RECT  7.38 6.30 7.74 6.66 ;
        RECT  4.14 5.22 4.50 5.58 ;
        RECT  1.98 6.30 2.34 6.66 ;
        LAYER metal2 ;
        RECT  7.26 5.10 7.86 5.70 ;
        RECT  4.02 5.10 4.62 5.70 ;
        RECT  4.02 5.16 7.86 5.64 ;
        RECT  7.26 6.18 7.86 6.78 ;
        RECT  1.86 6.18 2.46 6.78 ;
        RECT  1.86 6.24 7.86 6.72 ;
    END
END xor2_1

MACRO xor2_2
    CLASS CORE ;
    FOREIGN xor2_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.64 BY 15.12 ;
    SYMMETRY x y  ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.10 2.76 5.58 4.80 ;
        RECT  5.16 7.80 5.64 12.36 ;
        RECT  5.10 4.32 6.72 4.80 ;
        RECT  6.24 4.32 6.72 8.28 ;
        RECT  5.16 7.80 6.72 8.28 ;
        END
    END op
    PIN ip2
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal2 ;
        RECT  0.78 6.18 1.38 6.78 ;
        RECT  0.78 6.24 5.70 6.72 ;
        RECT  5.10 6.18 5.70 6.78 ;
        LAYER metal1 ;
        RECT  0.78 6.18 1.38 6.78 ;
        RECT  5.10 6.18 5.70 6.78 ;
        LAYER via ;
        RECT  0.90 6.30 1.26 6.66 ;
        RECT  5.22 6.30 5.58 6.66 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE analog ;
        PORT
        LAYER metal2 ;
        RECT  2.94 8.34 3.54 8.94 ;
        RECT  2.94 8.40 7.86 8.88 ;
        RECT  7.26 8.34 7.86 8.94 ;
        LAYER metal1 ;
        RECT  2.94 8.34 3.54 8.94 ;
        RECT  7.26 8.34 7.86 8.94 ;
        LAYER via ;
        RECT  3.06 8.46 3.42 8.82 ;
        RECT  7.38 8.46 7.74 8.82 ;
        END
    END ip1
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.42 0.00 0.90 4.26 ;
        RECT  3.42 0.00 3.90 3.96 ;
        RECT  6.84 0.00 7.32 3.96 ;
        RECT  0.00 0.00 8.64 1.32 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.42 9.24 0.90 15.12 ;
        RECT  3.42 10.14 3.90 15.12 ;
        RECT  6.84 9.30 7.32 15.12 ;
        RECT  0.00 13.80 8.64 15.12 ;
        END
    END vdd
    OBS
        LAYER metal1 ;
        RECT  7.26 5.10 7.86 5.70 ;
        RECT  7.26 7.26 7.86 7.86 ;
        RECT  2.46 9.30 2.94 12.36 ;
        RECT  2.46 9.30 4.56 9.78 ;
        RECT  4.08 4.32 4.56 9.78 ;
        RECT  4.02 4.32 4.62 5.70 ;
        RECT  2.46 4.32 4.62 4.80 ;
        RECT  2.46 2.76 2.94 4.80 ;
        RECT  1.38 8.40 1.86 12.36 ;
        RECT  1.38 8.40 2.40 8.88 ;
        RECT  1.92 5.16 2.40 8.88 ;
        RECT  1.86 7.26 2.46 7.86 ;
        RECT  1.38 5.16 2.40 5.64 ;
        RECT  1.38 2.76 1.86 5.64 ;
        LAYER via ;
        RECT  7.38 5.22 7.74 5.58 ;
        RECT  7.38 7.38 7.74 7.74 ;
        RECT  4.14 5.22 4.50 5.58 ;
        RECT  1.98 7.38 2.34 7.74 ;
        LAYER metal2 ;
        RECT  7.26 5.10 7.86 5.70 ;
        RECT  4.02 5.10 4.62 5.70 ;
        RECT  4.02 5.16 7.86 5.64 ;
        RECT  7.26 7.26 7.86 7.86 ;
        RECT  1.86 7.26 2.46 7.86 ;
        RECT  1.86 7.32 7.86 7.80 ;
    END
END xor2_2


MACRO padgnd
  CLASS  PAD ;
  FOREIGN padgnd 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 90.000 BY 300.000 ;
  SYMMETRY X Y R90  ;
  SITE IOSite ;
  PIN vddm1
    DIRECTION INOUT ;
    USE POWER ; SHAPE FEEDTHRU ;
    PORT
      LAYER metal1 ;
        RECT 0.000 0.000 0.480 100.320 ;
        RECT 89.520 0.000 90.000 100.320 ;
    END
  END vddm1
  PIN vdd1
    DIRECTION INOUT ;
    USE POWER ; SHAPE FEEDTHRU ;
    PORT
      LAYER metal2 ;
        RECT 0.000 135.120 0.480 209.040 ;
        RECT 89.520 135.120 90.000 209.040 ;
    END
  END vdd1
  PIN vdd2
    DIRECTION INOUT ;
    USE POWER ; SHAPE FEEDTHRU ;
    PORT
      LAYER metal2 ;
        RECT 0.000 78.120 0.480 100.320 ;
        RECT 89.520 78.120 90.000 100.320 ;
    END
  END vdd2
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 37.560 0.000 52.440 0.480 ;
    END
  END gnd
  PIN pad
    DIRECTION INPUT ;
    PORT
      LAYER metal5 ;
        RECT 9.000 228.000 81.000 300.000 ;
    END
  END pad
  PIN vss1
    DIRECTION INOUT ;
    USE GROUND ; SHAPE FEEDTHRU ;
    PORT
      LAYER metal2 ;
        RECT 0.000 108.720 0.480 130.920 ;
        RECT 89.520 108.720 90.000 130.920 ;
    END
  END vss1
  PIN vssm1
    DIRECTION INOUT ;
    USE GROUND ; SHAPE FEEDTHRU ;
    PORT
      LAYER metal1 ;
        RECT 0.000 108.720 0.480 209.040 ;
        RECT 89.520 108.720 90.000 209.040 ;
    END
  END vssm1
  PIN vss2
    DIRECTION INOUT ;
    USE GROUND ; SHAPE FEEDTHRU ;
    PORT
      LAYER metal2 ;
        RECT 0.000 0.000 0.480 73.920 ;
        RECT 89.520 0.000 90.000 73.920 ;
    END
  END vss2
  OBS 
      LAYER metal1 ;
        RECT 0.180 209.700 89.820 299.820 ;
        RECT 0.180 100.980 89.820 108.060 ;
        RECT 1.140 1.140 88.860 299.820 ;
        RECT 53.100 0.180 88.860 299.820 ;
        RECT 1.140 0.180 36.900 299.820 ;
      LAYER metal4 ;
        RECT 0.240 0.240 89.760 299.760 ;
      LAYER metal5 ;
        RECT 81.900 0.240 89.760 299.760 ;
        RECT 0.240 0.240 89.760 227.100 ;
        RECT 0.240 0.240 8.100 299.760 ;
      LAYER metal2 ;
        RECT 0.240 209.820 89.760 299.760 ;
        RECT 0.240 101.100 89.760 107.940 ;
        RECT 1.260 1.260 88.740 299.760 ;
        RECT 53.220 0.240 88.740 299.760 ;
        RECT 1.260 0.240 36.780 299.760 ;
      LAYER metal3 ;
        RECT 0.240 209.820 89.760 299.760 ;
        RECT 0.240 131.700 89.760 134.340 ;
        RECT 0.240 101.100 89.760 107.940 ;
        RECT 0.240 74.700 89.760 77.340 ;
        RECT 1.260 0.240 88.740 299.760 ;
  END 
END padgnd

MACRO padbidirhe_025
  CLASS  PAD ;
  FOREIGN padbidirhe_025 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 90.000 BY 300.000 ;
  SYMMETRY X Y R90  ;
  SITE IOSite ;
  PIN vddm1
    DIRECTION INOUT ;
    USE POWER ; SHAPE FEEDTHRU ;
    PORT
      LAYER metal1 ;
        RECT 0.000 0.000 0.480 100.320 ;
        RECT 89.520 0.000 90.000 100.320 ;
    END
  END vddm1
  PIN oeb
    DIRECTION INPUT ;
    PORT
      LAYER metal2 ;
        RECT 19.980 0.000 21.360 0.480 ;
    END
  END oeb
  PIN dib
    DIRECTION OUTPUT ;
    PORT
      LAYER metal2 ;
        RECT 63.360 0.000 64.680 0.480 ;
    END
  END dib
  PIN do
    DIRECTION INPUT ;
    PORT
      LAYER metal2 ;
        RECT 26.280 0.000 27.600 0.480 ;
    END
  END do
  PIN vdd1
    DIRECTION INOUT ;
    USE POWER ; SHAPE FEEDTHRU ;
    PORT
      LAYER metal2 ;
        RECT 0.000 135.120 0.480 209.040 ;
        RECT 89.520 135.120 90.000 209.040 ;
    END
  END vdd1
  PIN vdd2
    DIRECTION INOUT ;
    USE POWER ; SHAPE FEEDTHRU ;
    PORT
      LAYER metal2 ;
        RECT 0.000 78.120 0.480 100.320 ;
        RECT 89.520 78.120 90.000 100.320 ;
    END
  END vdd2
  PIN vss1
    DIRECTION INOUT ;
    USE GROUND ; SHAPE FEEDTHRU ;
    PORT
      LAYER metal2 ;
        RECT 0.000 108.720 0.480 130.920 ;
        RECT 89.520 108.720 90.000 130.920 ;
    END
  END vss1
  PIN pad
    DIRECTION INOUT ;
    PORT
      LAYER metal5 ;
        RECT 9.000 228.000 81.000 300.000 ;
    END
  END pad
  PIN vssm1
    DIRECTION INOUT ;
    USE GROUND ; SHAPE FEEDTHRU ;
    PORT
      LAYER metal1 ;
        RECT 0.000 108.720 0.480 209.040 ;
        RECT 89.520 108.720 90.000 209.040 ;
    END
  END vssm1
  PIN vss2
    DIRECTION INOUT ;
    USE GROUND ; SHAPE FEEDTHRU ;
    PORT
      LAYER metal2 ;
        RECT 0.000 0.000 0.480 73.920 ;
        RECT 89.520 0.000 90.000 73.920 ;
    END
  END vss2
  PIN di
    DIRECTION OUTPUT ;
    PORT
      LAYER metal2 ;
        RECT 66.000 0.000 67.320 0.480 ;
    END
  END di
  OBS 
      LAYER metal1 ;
        RECT 0.180 209.700 89.820 299.820 ;
        RECT 0.180 100.980 89.820 108.060 ;
        RECT 1.140 0.180 88.860 299.820 ;
      LAYER metal4 ;
        RECT 0.240 0.240 89.760 299.760 ;
      LAYER metal5 ;
        RECT 81.900 0.240 89.760 299.760 ;
        RECT 0.240 0.240 89.760 227.100 ;
        RECT 0.240 0.240 8.100 299.760 ;
      LAYER metal2 ;
        RECT 0.240 209.820 89.760 299.760 ;
        RECT 0.240 101.100 89.760 107.940 ;
        RECT 1.260 1.260 88.740 299.760 ;
        RECT 68.100 0.240 88.740 299.760 ;
        RECT 28.380 0.240 62.580 299.760 ;
        RECT 22.140 0.240 25.500 299.760 ;
        RECT 1.260 0.240 19.200 299.760 ;
      LAYER metal3 ;
        RECT 0.240 209.820 89.760 299.760 ;
        RECT 0.240 131.700 89.760 134.340 ;
        RECT 0.240 101.100 89.760 107.940 ;
        RECT 0.240 74.700 89.760 77.340 ;
        RECT 1.260 1.260 88.740 299.760 ;
        RECT 68.100 0.240 88.740 299.760 ;
        RECT 28.380 0.240 62.580 299.760 ;
        RECT 22.140 0.240 25.500 299.760 ;
        RECT 1.260 0.240 19.200 299.760 ;
  END 
END padbidirhe_025

MACRO padinc
  CLASS  PAD ;
  FOREIGN padinc 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 90.000 BY 300.000 ;
  SYMMETRY X Y R90  ;
  SITE IOSite ;
  PIN vddm1
    DIRECTION INOUT ;
    USE POWER ; SHAPE FEEDTHRU ;
    PORT
      LAYER metal1 ;
        RECT 0.000 0.000 0.480 100.320 ;
        RECT 89.520 0.000 90.000 100.320 ;
    END
  END vddm1
  PIN dib
    DIRECTION OUTPUT ;
    PORT
      LAYER metal2 ;
        RECT 63.360 0.000 64.680 0.480 ;
    END
  END dib
  PIN vdd1
    DIRECTION INOUT ;
    USE POWER ; SHAPE FEEDTHRU ;
    PORT
      LAYER metal2 ;
        RECT 0.000 135.120 0.480 209.040 ;
        RECT 89.520 135.120 90.000 209.040 ;
    END
  END vdd1
  PIN vdd2
    DIRECTION INOUT ;
    USE POWER ; SHAPE FEEDTHRU ;
    PORT
      LAYER metal2 ;
        RECT 0.000 78.120 0.480 100.320 ;
        RECT 89.520 78.120 90.000 100.320 ;
    END
  END vdd2
  PIN vss1
    DIRECTION INOUT ;
    USE GROUND ; SHAPE FEEDTHRU ;
    PORT
      LAYER metal2 ;
        RECT 0.000 108.720 0.480 130.920 ;
        RECT 89.520 108.720 90.000 130.920 ;
    END
  END vss1
  PIN pad
    DIRECTION INPUT ;
    PORT
      LAYER metal5 ;
        RECT 9.000 228.000 81.000 300.000 ;
    END
  END pad
  PIN vssm1
    DIRECTION INOUT ;
    USE GROUND ; SHAPE FEEDTHRU ;
    PORT
      LAYER metal1 ;
        RECT 0.000 108.720 0.480 209.040 ;
        RECT 89.520 108.720 90.000 209.040 ;
    END
  END vssm1
  PIN vss2
    DIRECTION INOUT ;
    USE GROUND ; SHAPE FEEDTHRU ;
    PORT
      LAYER metal2 ;
        RECT 0.000 0.000 0.480 73.920 ;
        RECT 89.520 0.000 90.000 73.920 ;
    END
  END vss2
  PIN di
    DIRECTION OUTPUT ;
    PORT
      LAYER metal2 ;
        RECT 66.000 0.000 67.320 0.480 ;
    END
  END di
  OBS 
      LAYER metal1 ;
        RECT 0.180 209.700 89.820 299.820 ;
        RECT 0.180 100.980 89.820 108.060 ;
        RECT 1.140 0.180 88.860 299.820 ;
      LAYER metal4 ;
        RECT 0.240 0.240 89.760 299.760 ;
      LAYER metal5 ;
        RECT 81.900 0.240 89.760 299.760 ;
        RECT 0.240 0.240 89.760 227.100 ;
        RECT 0.240 0.240 8.100 299.760 ;
      LAYER metal2 ;
        RECT 0.240 209.820 89.760 299.760 ;
        RECT 0.240 101.100 89.760 107.940 ;
        RECT 1.260 1.260 88.740 299.760 ;
        RECT 68.100 0.240 88.740 299.760 ;
        RECT 1.260 0.240 62.580 299.760 ;
      LAYER metal3 ;
        RECT 0.240 209.820 89.760 299.760 ;
        RECT 0.240 131.700 89.760 134.340 ;
        RECT 0.240 101.100 89.760 107.940 ;
        RECT 0.240 74.700 89.760 77.340 ;
        RECT 1.260 1.260 88.740 299.760 ;
        RECT 68.100 0.240 88.740 299.760 ;
        RECT 1.260 0.240 62.580 299.760 ;
  END 
END padinc

MACRO padio
  CLASS  PAD ;
  FOREIGN padio 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 90.000 BY 300.000 ;
  SYMMETRY X Y R90  ;
  SITE IOSite ;
  PIN vddm1
    DIRECTION INOUT ;
    USE POWER ; SHAPE FEEDTHRU ;
    PORT
      LAYER metal1 ;
        RECT 0.000 0.000 0.480 100.320 ;
        RECT 89.520 0.000 90.000 100.320 ;
    END
  END vddm1
  PIN data
    DIRECTION INOUT ;
    PORT
      LAYER metal2 ;
        RECT 37.560 0.000 52.440 0.480 ;
    END
  END data
  PIN vdd1
    DIRECTION INOUT ;
    USE POWER ; SHAPE FEEDTHRU ;
    PORT
      LAYER metal2 ;
        RECT 0.000 135.120 0.480 209.040 ;
        RECT 89.520 135.120 90.000 209.040 ;
    END
  END vdd1
  PIN vdd2
    DIRECTION INOUT ;
    USE POWER ; SHAPE FEEDTHRU ;
    PORT
      LAYER metal2 ;
        RECT 0.000 78.120 0.480 100.320 ;
        RECT 89.520 78.120 90.000 100.320 ;
    END
  END vdd2
  PIN vss1
    DIRECTION INOUT ;
    USE GROUND ; SHAPE FEEDTHRU ;
    PORT
      LAYER metal2 ;
        RECT 0.000 108.720 0.480 130.920 ;
        RECT 89.520 108.720 90.000 130.920 ;
    END
  END vss1
  PIN pad
    DIRECTION INOUT ;
    PORT
      LAYER metal5 ;
        RECT 9.000 228.000 81.000 300.000 ;
    END
  END pad
  PIN vssm1
    DIRECTION INOUT ;
    USE GROUND ; SHAPE FEEDTHRU ;
    PORT
      LAYER metal1 ;
        RECT 0.000 108.720 0.480 209.040 ;
        RECT 89.520 108.720 90.000 209.040 ;
    END
  END vssm1
  PIN vss2
    DIRECTION INOUT ;
    USE GROUND ; SHAPE FEEDTHRU ;
    PORT
      LAYER metal2 ;
        RECT 0.000 0.000 0.480 73.920 ;
        RECT 89.520 0.000 90.000 73.920 ;
    END
  END vss2
  OBS 
      LAYER metal1 ;
        RECT 0.180 209.700 89.820 299.820 ;
        RECT 0.180 100.980 89.820 108.060 ;
        RECT 1.140 0.180 88.860 299.820 ;
      LAYER metal4 ;
        RECT 0.240 0.240 89.760 299.760 ;
      LAYER metal5 ;
        RECT 81.900 0.240 89.760 299.760 ;
        RECT 0.240 0.240 89.760 227.100 ;
        RECT 0.240 0.240 8.100 299.760 ;
      LAYER metal2 ;
        RECT 0.240 209.820 89.760 299.760 ;
        RECT 0.240 101.100 89.760 107.940 ;
        RECT 1.260 1.260 88.740 299.760 ;
        RECT 53.220 0.240 88.740 299.760 ;
        RECT 1.260 0.240 36.780 299.760 ;
      LAYER metal3 ;
        RECT 0.240 209.820 89.760 299.760 ;
        RECT 0.240 131.700 89.760 134.340 ;
        RECT 0.240 101.100 89.760 107.940 ;
        RECT 0.240 74.700 89.760 77.340 ;
        RECT 1.260 1.260 88.740 299.760 ;
        RECT 53.220 0.240 88.740 299.760 ;
        RECT 1.260 0.240 36.780 299.760 ;
  END 
END padio

MACRO padlesscorner
  CLASS  ENDCAP TOPLEFT ;
  FOREIGN padlesscorner 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 300.000 ;
  SYMMETRY X Y R90  ;
  SITE CornerSite ;
  PIN vddm1
    DIRECTION INOUT ;
    USE POWER ; SHAPE FEEDTHRU ;
    PORT
      LAYER metal1 ;
        RECT 199.680 0.000 300.000 0.480 ;
        RECT 299.520 0.000 300.000 100.320 ;
    END
  END vddm1
  PIN vdd1
    DIRECTION INOUT ;
    USE POWER ; SHAPE FEEDTHRU ;
    PORT
      LAYER metal2 ;
        RECT 90.960 0.000 164.880 0.480 ;
        RECT 299.520 135.120 300.000 209.040 ;
    END
  END vdd1
  PIN vdd2
    DIRECTION INOUT ;
    USE POWER ; SHAPE FEEDTHRU ;
    PORT
      LAYER metal2 ;
        RECT 199.680 0.000 221.880 0.480 ;
        RECT 299.520 78.120 300.000 100.320 ;
    END
  END vdd2
  PIN vss1
    DIRECTION INOUT ;
    USE GROUND ; SHAPE FEEDTHRU ;
    PORT
      LAYER metal2 ;
        RECT 169.080 0.000 191.280 0.480 ;
        RECT 299.520 108.720 300.000 130.920 ;
    END
  END vss1
  PIN vssm1
    DIRECTION INOUT ;
    USE GROUND ; SHAPE FEEDTHRU ;
    PORT
      LAYER metal1 ;
        RECT 90.960 0.000 191.280 0.480 ;
        RECT 299.520 108.720 300.000 209.040 ;
    END
  END vssm1
  PIN vss2
    DIRECTION INOUT ;
    USE GROUND ; SHAPE FEEDTHRU ;
    PORT
      LAYER metal2 ;
        RECT 226.080 0.000 300.000 0.480 ;
        RECT 299.520 0.000 300.000 73.920 ;
    END
  END vss2
  OBS 
      LAYER metal1 ;
        RECT 0.180 209.700 299.820 299.820 ;
        RECT 0.180 100.980 299.820 108.060 ;
        RECT 0.180 1.140 298.860 299.820 ;
        RECT 191.940 0.180 199.020 299.820 ;
        RECT 0.180 0.180 90.300 299.820 ;
      LAYER metal4 ;
        RECT 0.240 0.240 299.760 299.760 ;
      LAYER metal5 ;
        RECT 0.240 0.240 299.760 299.760 ;
      LAYER metal2 ;
        RECT 0.240 209.820 299.760 299.760 ;
        RECT 0.240 101.100 299.760 107.940 ;
        RECT 0.240 1.260 298.740 299.760 ;
        RECT 192.060 0.240 198.900 299.760 ;
        RECT 0.240 0.240 90.180 299.760 ;
      LAYER metal3 ;
        RECT 0.240 209.820 299.760 299.760 ;
        RECT 0.240 131.700 299.760 134.340 ;
        RECT 0.240 101.100 299.760 107.940 ;
        RECT 0.240 74.700 299.760 77.340 ;
        RECT 0.240 1.260 298.740 299.760 ;
        RECT 222.660 0.240 225.300 299.760 ;
        RECT 192.060 0.240 198.900 299.760 ;
        RECT 165.660 0.240 168.300 299.760 ;
        RECT 0.240 0.240 90.180 299.760 ;
  END 
END padlesscorner

MACRO padout
  CLASS  PAD ;
  FOREIGN padout 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 90.000 BY 300.000 ;
  SYMMETRY X Y R90  ;
  SITE IOSite ;
  PIN vddm1
    DIRECTION INOUT ;
    USE POWER ; SHAPE FEEDTHRU ;
    PORT
      LAYER metal1 ;
        RECT 0.000 0.000 0.480 100.320 ;
        RECT 89.520 0.000 90.000 100.320 ;
    END
  END vddm1
  PIN dib
    DIRECTION OUTPUT ;
    PORT
      LAYER metal2 ;
        RECT 63.360 0.000 64.680 0.480 ;
    END
  END dib
  PIN do
    DIRECTION INPUT ;
    PORT
      LAYER metal2 ;
        RECT 26.280 0.000 27.600 0.480 ;
    END
  END do
  PIN vdd1
    DIRECTION INOUT ;
    USE POWER ; SHAPE FEEDTHRU ;
    PORT
      LAYER metal2 ;
        RECT 0.000 135.120 0.480 209.040 ;
        RECT 89.520 135.120 90.000 209.040 ;
    END
  END vdd1
  PIN vdd2
    DIRECTION INOUT ;
    USE POWER ; SHAPE FEEDTHRU ;
    PORT
      LAYER metal2 ;
        RECT 0.000 78.120 0.480 100.320 ;
        RECT 89.520 78.120 90.000 100.320 ;
    END
  END vdd2
  PIN vss1
    DIRECTION INOUT ;
    USE GROUND ; SHAPE FEEDTHRU ;
    PORT
      LAYER metal2 ;
        RECT 0.000 108.720 0.480 130.920 ;
        RECT 89.520 108.720 90.000 130.920 ;
    END
  END vss1
  PIN pad
    DIRECTION OUTPUT ;
    PORT
      LAYER metal5 ;
        RECT 9.000 228.000 81.000 300.000 ;
    END
  END pad
  PIN vssm1
    DIRECTION INOUT ;
    USE GROUND ; SHAPE FEEDTHRU ;
    PORT
      LAYER metal1 ;
        RECT 0.000 108.720 0.480 209.040 ;
        RECT 89.520 108.720 90.000 209.040 ;
    END
  END vssm1
  PIN vss2
    DIRECTION INOUT ;
    USE GROUND ; SHAPE FEEDTHRU ;
    PORT
      LAYER metal2 ;
        RECT 0.000 0.000 0.480 73.920 ;
        RECT 89.520 0.000 90.000 73.920 ;
    END
  END vss2
  PIN di
    DIRECTION OUTPUT ;
    PORT
      LAYER metal2 ;
        RECT 66.000 0.000 67.320 0.480 ;
    END
  END di
  OBS 
      LAYER metal1 ;
        RECT 0.180 209.700 89.820 299.820 ;
        RECT 0.180 100.980 89.820 108.060 ;
        RECT 1.140 0.180 88.860 299.820 ;
      LAYER metal4 ;
        RECT 0.240 0.240 89.760 299.760 ;
      LAYER metal5 ;
        RECT 81.900 0.240 89.760 299.760 ;
        RECT 0.240 0.240 89.760 227.100 ;
        RECT 0.240 0.240 8.100 299.760 ;
      LAYER metal2 ;
        RECT 0.240 209.820 89.760 299.760 ;
        RECT 0.240 101.100 89.760 107.940 ;
        RECT 1.260 1.260 88.740 299.760 ;
        RECT 68.100 0.240 88.740 299.760 ;
        RECT 28.380 0.240 62.580 299.760 ;
        RECT 1.260 0.240 25.500 299.760 ;
      LAYER metal3 ;
        RECT 0.240 209.820 89.760 299.760 ;
        RECT 0.240 131.700 89.760 134.340 ;
        RECT 0.240 101.100 89.760 107.940 ;
        RECT 0.240 74.700 89.760 77.340 ;
        RECT 1.260 1.260 88.740 299.760 ;
        RECT 68.100 0.240 88.740 299.760 ;
        RECT 28.380 0.240 62.580 299.760 ;
        RECT 1.260 0.240 25.500 299.760 ;
  END 
END padout

MACRO padvdd
  CLASS  PAD ;
  FOREIGN padvdd 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 90.000 BY 300.000 ;
  SYMMETRY X Y R90  ;
  SITE IOSite ;
  PIN vddm1
    DIRECTION INOUT ;
    USE POWER ; SHAPE FEEDTHRU ;
    PORT
      LAYER metal1 ;
        RECT 0.000 0.000 0.480 100.320 ;
        RECT 89.520 0.000 90.000 100.320 ;
    END
  END vddm1
  PIN vdd1
    DIRECTION INOUT ;
    USE POWER ; SHAPE FEEDTHRU ;
    PORT
      LAYER metal2 ;
        RECT 0.000 135.120 0.480 209.040 ;
        RECT 89.520 135.120 90.000 209.040 ;
    END
  END vdd1
  PIN vdd2
    DIRECTION INOUT ;
    USE POWER ; SHAPE FEEDTHRU ;
    PORT
      LAYER metal2 ;
        RECT 0.000 78.120 0.480 100.320 ;
        RECT 89.520 78.120 90.000 100.320 ;
    END
  END vdd2
  PIN vss1
    DIRECTION INOUT ;
    USE GROUND ; SHAPE FEEDTHRU ;
    PORT
      LAYER metal2 ;
        RECT 0.000 108.720 0.480 130.920 ;
        RECT 89.520 108.720 90.000 130.920 ;
    END
  END vss1
  PIN pad
    DIRECTION INPUT ;
    PORT
      LAYER metal5 ;
        RECT 9.000 228.000 81.000 300.000 ;
    END
  END pad
  PIN vssm1
    DIRECTION INOUT ;
    USE GROUND ; SHAPE FEEDTHRU ;
    PORT
      LAYER metal1 ;
        RECT 0.000 108.720 0.480 209.040 ;
        RECT 89.520 108.720 90.000 209.040 ;
    END
  END vssm1
  PIN vss2
    DIRECTION INOUT ;
    USE GROUND ; SHAPE FEEDTHRU ;
    PORT
      LAYER metal2 ;
        RECT 0.000 0.000 0.480 73.920 ;
        RECT 89.520 0.000 90.000 73.920 ;
    END
  END vss2
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 37.560 0.000 52.440 0.480 ;
    END
  END vdd
  OBS 
      LAYER metal1 ;
        RECT 0.180 209.700 89.820 299.820 ;
        RECT 0.180 100.980 89.820 108.060 ;
        RECT 1.140 1.140 88.860 299.820 ;
        RECT 53.100 0.180 88.860 299.820 ;
        RECT 1.140 0.180 36.900 299.820 ;
      LAYER metal4 ;
        RECT 0.240 0.240 89.760 299.760 ;
      LAYER metal5 ;
        RECT 81.900 0.240 89.760 299.760 ;
        RECT 0.240 0.240 89.760 227.100 ;
        RECT 0.240 0.240 8.100 299.760 ;
      LAYER metal2 ;
        RECT 0.240 209.820 89.760 299.760 ;
        RECT 0.240 101.100 89.760 107.940 ;
        RECT 1.260 1.260 88.740 299.760 ;
        RECT 53.220 0.240 88.740 299.760 ;
        RECT 1.260 0.240 36.780 299.760 ;
      LAYER metal3 ;
        RECT 0.240 209.820 89.760 299.760 ;
        RECT 0.240 131.700 89.760 134.340 ;
        RECT 0.240 101.100 89.760 107.940 ;
        RECT 0.240 74.700 89.760 77.340 ;
        RECT 1.260 0.240 88.740 299.760 ;
  END 
END padvdd

MACRO padnoconnect
  CLASS  PAD ;
  FOREIGN padnoconnect 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 90.000 BY 300.000 ;
  SYMMETRY X Y R90  ;
  SITE IOSite ;
  PIN vddm1
    DIRECTION INOUT ;
    USE POWER ; SHAPE FEEDTHRU ;
    PORT
      LAYER metal1 ;
        RECT 0.000 0.000 0.480 100.320 ;
        RECT 89.520 0.000 90.000 100.320 ;
    END
  END vddm1
  PIN vdd1
    DIRECTION INOUT ;
    USE POWER ; SHAPE FEEDTHRU ;
    PORT
      LAYER metal2 ;
        RECT 0.000 135.120 0.480 209.040 ;
        RECT 89.520 135.120 90.000 209.040 ;
    END
  END vdd1
  PIN vdd2
    DIRECTION INOUT ;
    USE POWER ; SHAPE FEEDTHRU ;
    PORT
      LAYER metal2 ;
        RECT 0.000 78.120 0.480 100.320 ;
        RECT 89.520 78.120 90.000 100.320 ;
    END
  END vdd2
  PIN vss1
    DIRECTION INOUT ;
    USE GROUND ; SHAPE FEEDTHRU ;
    PORT
      LAYER metal2 ;
        RECT 0.000 108.720 0.480 130.920 ;
        RECT 89.520 108.720 90.000 130.920 ;
    END
  END vss1
  PIN pad
    DIRECTION INPUT ;
    PORT
      LAYER metal5 ;
        RECT 9.000 228.000 81.000 300.000 ;
    END
  END pad
  PIN vssm1
    DIRECTION INOUT ;
    USE GROUND ; SHAPE FEEDTHRU ;
    PORT
      LAYER metal1 ;
        RECT 0.000 108.720 0.480 209.040 ;
        RECT 89.520 108.720 90.000 209.040 ;
    END
  END vssm1
  PIN vss2
    DIRECTION INOUT ;
    USE GROUND ; SHAPE FEEDTHRU ;
    PORT
      LAYER metal2 ;
        RECT 0.000 0.000 0.480 73.920 ;
        RECT 89.520 0.000 90.000 73.920 ;
    END
  END vss2
  OBS 
      LAYER metal1 ;
        RECT 0.180 209.700 89.820 299.820 ;
        RECT 0.180 100.980 89.820 108.060 ;
        RECT 1.140 0.180 88.860 299.820 ;
      LAYER metal4 ;
        RECT 0.240 0.240 89.760 299.760 ;
      LAYER metal5 ;
        RECT 81.900 0.240 89.760 299.760 ;
        RECT 0.240 0.240 89.760 227.100 ;
        RECT 0.240 0.240 8.100 299.760 ;
      LAYER metal2 ;
        RECT 0.240 209.820 89.760 299.760 ;
        RECT 0.240 101.100 89.760 107.940 ;
        RECT 1.260 0.240 88.740 299.760 ;
      LAYER metal3 ;
        RECT 0.240 209.820 89.760 299.760 ;
        RECT 0.240 131.700 89.760 134.340 ;
        RECT 0.240 101.100 89.760 107.940 ;
        RECT 0.240 74.700 89.760 77.340 ;
        RECT 1.260 0.240 88.740 299.760 ;
  END 
END padnoconnect

MACRO padlessspacer
  CLASS  PAD ;
  FOREIGN padlessspacer 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 90.000 BY 300.000 ;
  SYMMETRY X Y R90  ;
  SITE IOSite ;
  PIN vddm1
    DIRECTION INOUT ;
    USE POWER ; SHAPE FEEDTHRU ;
    PORT
      LAYER metal1 ;
        RECT 0.000 0.000 0.480 100.320 ;
        RECT 89.520 0.000 90.000 100.320 ;
    END
  END vddm1
  PIN vdd1
    DIRECTION INOUT ;
    USE POWER ; SHAPE FEEDTHRU ;
    PORT
      LAYER metal2 ;
        RECT 0.000 135.120 0.480 209.040 ;
        RECT 89.520 135.120 90.000 209.040 ;
    END
  END vdd1
  PIN vdd2
    DIRECTION INOUT ;
    USE POWER ; SHAPE FEEDTHRU ;
    PORT
      LAYER metal2 ;
        RECT 0.000 78.120 0.480 100.320 ;
        RECT 89.520 78.120 90.000 100.320 ;
    END
  END vdd2
  PIN vss1
    DIRECTION INOUT ;
    USE GROUND ; SHAPE FEEDTHRU ;
    PORT
      LAYER metal2 ;
        RECT 0.000 108.720 0.480 130.920 ;
        RECT 89.520 108.720 90.000 130.920 ;
    END
  END vss1
  PIN vssm1
    DIRECTION INOUT ;
    USE GROUND ; SHAPE FEEDTHRU ;
    PORT
      LAYER metal1 ;
        RECT 0.000 108.720 0.480 209.040 ;
        RECT 89.520 108.720 90.000 209.040 ;
    END
  END vssm1
  PIN vss2
    DIRECTION INOUT ;
    USE GROUND ; SHAPE FEEDTHRU ;
    PORT
      LAYER metal2 ;
        RECT 0.000 0.000 0.480 73.920 ;
        RECT 89.520 0.000 90.000 73.920 ;
    END
  END vss2
  OBS 
      LAYER metal1 ;
        RECT 0.180 209.700 89.820 299.820 ;
        RECT 0.180 100.980 89.820 108.060 ;
        RECT 1.140 0.180 88.860 299.820 ;
      LAYER metal4 ;
        RECT 0.240 0.240 89.760 299.760 ;
      LAYER metal5 ;
        RECT 0.240 0.240 89.760 299.760 ;
      LAYER metal2 ;
        RECT 0.240 209.820 89.760 299.760 ;
        RECT 0.240 101.100 89.760 107.940 ;
        RECT 1.260 0.240 88.740 299.760 ;
      LAYER metal3 ;
        RECT 0.240 209.820 89.760 299.760 ;
        RECT 0.240 131.700 89.760 134.340 ;
        RECT 0.240 101.100 89.760 107.940 ;
        RECT 0.240 74.700 89.760 77.340 ;
        RECT 1.260 0.240 88.740 299.760 ;
  END 
END padlessspacer

END LIBRARY
