// ECE 425 MP2: Verilog RTL for Am2901 controller
// Rev 2/17/08

module controller(
	i,					// opcode (add your decoded signals)
	a,b,select_a_hi,select_b_hi,		// decoding of register addresses
	f,c,p,g_lo,p_lo,ovr,z,			// generation of ALU outputs
	y_tri,y_data,oe,			// tristate control of y bus
	ram0,ram3,		// tristate control of RAM shifter
	q0,q3,q0_data,q3_data,			// tristate control of Q shifter
	reg_wr,      //write_en for RAM. 
	r_sel, s_sel, func_sel, //Select signals to choose what we want ALU sources and function to be.
	y_sel, f_sel, q_sel, //Select signals for output and Q reg and RAM.
	zero, q_en,	//Zero = 0, q_en is for when we write to Q reg
	inv_s, inv_r,	//Inverts our s,r signals if set
	q_master_en, q_slave_en, iq_master_en, iq_slave_en, ireg_wr,
	reg_a_wr, ireg_a_wr, reg_b_wr, ireg_b_wr,
	cp
);

 // define I/O for synthesized control
input [8:0] i;
input [3:0] a, b;
output [15:0] select_a_hi, select_b_hi;
input [3:0] f, c, p;
output g_lo, p_lo, ovr, z;
inout [3:0] y_tri;
input [3:0] y_data;
input oe;
inout ram0, ram3, q0, q3;
input q0_data, q3_data;
output reg_wr;      //write_en for RAM. 
output reg [1:0] r_sel, s_sel, f_sel, q_sel; 
output [2:0] func_sel; //Select signals to choose what we want ALU sources and function to be.
output y_sel; //Select signals for output and Q reg and RAM.
output zero, q_en;	//Zero = 0, q_en is for when we write to Q reg
output inv_s, inv_r;
output q_master_en, q_slave_en, iq_master_en, iq_slave_en, ireg_wr;
input cp;
output reg_a_wr, ireg_a_wr, reg_b_wr, ireg_b_wr;

 // named internal wires carry reusable subexpressions
wire shift_left, shift_right;

 // "assign" statements give us algebraic expressions
assign select_a_hi = (16'h0001 << a);
assign select_b_hi = (16'h0001 << b);
assign shift_left = i[8] & i[7];
assign shift_right = i[8] & ~ i[7];

 // simpler functionality is better implemented directly in logic gates
buf calcg(	g_lo,	~c[3] ); // glitchy with lookahead carry propagation, but shouldn't matter for us :v)
nand calcp(	p_lo,	p[3], p[2], p[1], p[0] );
xor calcovr(	ovr,	c[3], c[2] );
nor calczero(	z,	f[3], f[2], f[1], f[0] );

bufif1 drvy3(	y_tri[3],y_data[3], oe );
bufif1 drvy2(	y_tri[2],y_data[2], oe );
bufif1 drvy1(	y_tri[1],y_data[1], oe );
bufif1 drvy0(	y_tri[0],y_data[0], oe );
bufif1 drvraml( ram3,	f[3], shift_left );
bufif1 drvramr( ram0,	f[0], shift_right );
bufif1 drvqshl( q3,	q3_data, shift_left );
bufif1 drvqshr( q0,	q0_data, shift_right );


 // add your control signals here...
always @(*) //Combinational
	begin
		r_sel = 2'b00; //Default
		s_sel = 2'b00; //Default
		f_sel = 2'b00; //Default
		q_sel = 2'b00; //Default
		if ( i[2] & (i[1] | i[0]) ) //r_sel = 0
			r_sel = 2'b00;
		else if ( (~i[2] & ~i[1]) ) //r_sel = 1
			r_sel = 2'b01;
		else if ( (~i[2] & i[1]) | (i[2] & ~i[1] & ~i[0]) ) //r_sel = 2
			r_sel = 2'b10;
		else
			r_sel = 2'b00;
		//s_sel
		if (i[2] & ~i[1])
			s_sel = 2'b00; 
		else if (~i[2] & i[0])
			s_sel = 2'b01;
		else if ( ~i[0] & ((i[2] & i[1]) | ~i[2]))
			s_sel = 2'b10;
		else if (i[2] & i[1] & i[0])
			s_sel = 2'b11;
		else
			s_sel = 2'b00;
		//f_sel
		if (i[8] & ~i[7])
			f_sel = 2'b00;
		else if (~i[8] & i[7])
			f_sel = 2'b01;
		else if (i[8] & i[7])
			f_sel = 2'b10;
		else
			f_sel = 2'b00; 
		//q_sel
		if (i[8] & ~i[7] & ~i[6])
			q_sel = 2'b00; //(Q >> 1) --> 0Q. Shift right
		else if (~i[8] & ~i[7] & ~i[6])
			q_sel = 2'b01; //F --> Q. Load
		else if (i[8] & i[7] & ~i[6])
			q_sel = 2'b10; //(Q << 1) --> Q. Shift left.
		else
			q_sel = 2'b00; 
	end
assign func_sel = {i[5], i[4], i[3]};
assign y_sel = ~(~i[8] & i[7] & ~i[6]); //Select signals for output and Q reg and RAM.
assign zero = 1'b0;
assign q_master_en = ((~i[8] & ~i[7] & ~i[6]) | (i[8] & ~i[7] & ~i[6]) | (i[8] & i[7] & ~i[6])) & ~cp;	
assign iq_master_en = ~q_master_en;

assign inv_s = (~i[5] & ~i[4] & ~i[3]) | (~i[5] & ~i[4] & i[3]) | (i[5] & i[4]); //~5~4~3=ADD, ~5~43=SUBR, 54=XOR,XNOR
assign inv_r = (~i[5] & ~i[4] & ~i[3]) | (~i[5] & i[4] & ~i[3]) | (i[5] & i[4]) | (i[5] & ~i[4] & i[3]) /*| (~i[5] & ~i[4] & i[3])*/;
assign reg_wr = (i[8] | i[7]) & ~cp;
assign ireg_wr = ~reg_wr;

assign q_slave_en = ((~i[8] & ~i[7] & ~i[6]) | (i[8] & ~i[7] & ~i[6]) | (i[8] & i[7] & ~i[6])) & cp;
assign iq_slave_en = ~q_slave_en;
assign reg_a_wr = cp;
assign ireg_a_wr = ~reg_a_wr;
assign reg_b_wr = cp;
assign ireg_b_wr = ~reg_b_wr;
endmodule

